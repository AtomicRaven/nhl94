GST@�                                                            \     �                                                ����      �  ��  �         ����e ����J�������ĸ����������        Fi     #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    
 �j,� B ��
  >�                                                                              ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������=o  0  4g  1                      �                         �  �  �  �                  �  
          8 �����������������������������������������������������������������������������                                ,x  q   n  ��   @  #   �   �                                                                                '       )n)n1n  
�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    Lb�WLCTs���h��T|7�AQ�QAlJQ|��)�t@ T0 k� �0 �4 %e1d  3Ab5p�  ��(    � 9 �Lb�WLCTs�� h��T|7�AQ�QAlJQt ��)�x@ T0 k� �, �0 %e1d  3Ab5p�  ��(    � 9 �Lb�WLC Ts�� g��T|7�AQ�QAlJQp ��)�x@ T0 k� �( �, %e1d  3Ab5p�  ��(    � 9 �Lb�WLC Ts��g��T|7�AQ�QAhJQl ��)�|@ T0 k� �  �$ %e1d  3Ab5p�  ��(    � 9 �Lb�WLC Ts��g��T|7�AQ�RAhJQd ��)�|@ T0 k� ���#�%e1d  3Ab5p�  ��(    � 9 �Lb�WLC Ts��g��T|7�AQ�RAhJQ` ��)�|@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �Lb�WLB�Ts��g��T|7�AQ�RAhJQ\ ��)À@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �Lb�WLB�Ts��f��T|7�AQ�RAhJQX ��)À@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �Lb�WLB�Ts��f��T|7�AQ�RAhJQP ��)À@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �Lb�VLB�Ts��f¸T|7�AQ�RAhJQO���)Ä@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �Lb�VLB�Ts��f¸T|7�AQ�RAhJQK���)Ä@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �Lb�VLB�Ts��f¸T|7�AQ�RAhJQG���)Ä@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �Lb�VLB�Ts��f¸T|7�AQ�RAhJQC���)È@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �Lb�VLB�Ts��f¸T|7�AQ�RAhJQ?���*È@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �Lb�VLB�Ts��f¸T|7�AQ�RAhJQ;���*Ì@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�ULB�Ts��f¸T|7�AQ�RAhJQ3���*Ì@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�ULB�Ts��f¸T|7�AQ�RAhJQ/���*Ì@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�ULB�Ts��f¸T|7�AQ�RAhJQ+���*Ð@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�ULB�Ts��f¸T|7�AQ�RAhJQ'���*Ð@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�ULB�Ts��f¸T|7�AQ�RAhJQ#���*Ð@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�ULB�Ts��f¸T|7�AQ�RAhJQ���*Ð@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�ULB�Ts��f¸T|7�AQ�RAhJQ���*Ô@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�TLB�Ts��f¸T|7�AQ�RAdJQ���*Ô@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�TLB�To��f¸T|7�AQ�RAdJQ���*Ô@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �LR�TLB�To��f¸T|7�AQ�RAdJQ���*Ø@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�RAdJQ���*Ø@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�RAdJQ���*Ø@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�RAdJQ���*Ø@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�RAdJQ���*Ü@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�RAdJP����*Ü@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�RAdJP����*Ü@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�RAdJP����*à@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�RAdJP����*à@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�RAdJP����*à@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�SAdJP����*à@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TLB�To��f¸T|7�AQ�SAdJP����*ä@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TL2�To��f¸T|7�AQ�SAdJP����*ä@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TL2�To��f¸T|7�AQ�SAdJP����*ä@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TL2�To��f¸T|7�AQ�SAdJP����*ä@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TL2�To��f¸T|7�AQ�SAdJP����*ä@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �A��TL2�o��f¸T|7�AQ�SAdJP����*è@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �A��TL2�o��f¸T|7�AQ�SAdJP����*è@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �A��TD2�o��f¸T|7�AQ|SAdJP����*è@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �A��TD2�o��f¸T|7�AQ|SAdJP����*è@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �AR�TD2�o��f¸T|7�AQ|SAdJP����*ì@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �AR�TD2�o��f¸T|7�AQ|SAdJP����*ì@ T0 k� ������%e1d  3Ab5p�  ��(    � 9 �AR�TD2�o��f¸T|7�AQ|SAdIP����*ì@ T0 k� �����%e1d  3Ab5p�  ��(    � 9 �AR�TD��o��f¸T|7�AQ|SAdIP����*ì@ T0 k� �{���%e1d  3Ab5p�  ��(    � 9 �AR�TD��o��f¸T|7�AQ|SAdIP����*ì@ T0 k� �{���%e1d  3Ab5p�  ��(   � 9 �AR�TD��o��f¸T|7�AQ|SAdIP����*ð@ T0 k� �w��{�%e1d  3Ab5p�  ��(    � 9 �AR�TD��o��f��T|7�AQ|SAdIP����*ð@ T0 k� �s��w�%e1d  3Ab5p�  ��(    � 9 �AR�TD��o��f��T|7�AQ|SA`IP����*ð@ T0 k� �s��w�%e1d  3Ab5p�  ��(    � 9 �AR�TD��o�3f��T|7�AQ|SA`IP����+ð@ T0 k� �o��s�%e1d  3Ab5p�  ��(    � 9 �AR�TD�� o�3f��T|7�AQ|SA`IP����+ð@ T0 k� �o��s�%e1d  3Ab5p�  ��(    � 9 �AR�TD�� $o�3f��T|7�AQ|SA`IP����+ô@ T0 k� �k��o�%e1d  3Ab5p�  ��(    � 9 �AR�TD�� $o�3f��T|7�AQ|SA`IP����+ô@ T0 k� �g��k�%e1d  3Ab5p�  ��(    � 9 �A�TD�� $o�3f b�T|7�AQ|SA`IP����+ô@ T0 k� �g��k�%e1d  3Ab5p�  ��(   � 9 �A�TD��!$o�3f b�T|7�AQ|SA`IP����+ô@ T0 k� �c��g�%e1d  3Ab5p�  ��(    � 9 �A�TD��!$o�3f b�T|7�AQxSA`IP����,ô@ T0 k� �c��g�%e1d  3Ab5p�  ��(    � 9 �A�TD��"$o�3f b�T|7�AQxSA`IP����,ô@ T0 k� �_��c�%e1d  3Ab5p�  ��(    � 9 �A�TD��"$o�3f b�T|7�AQxSA`IP����,ø@ T0 k� �_��c�%e1d  3Ab5p�  ��(    � 9 �A�TD��#$o�3f��T|7�AQxSA`IP����,ø@ T0 k� �[��_�%e1d  3Ab5p�  ��(    � 9 �A�TD��#$o�3f��T|7�AQxSA`IP����,ø@ T0 k� �[��_�%e1d  3Ab5p�  ��(    � 9 �A�TD��$$o�3f��T|7�AQxSA`IP����,ø@ T0 k� �W��[�%e1d  3Ab5p�  ��(    � 9 �A�TD��%$o�3f��T|7�AQxSA`IP����-ø@ T0 k� �W��[�%e1d  3Ab5p�  ��(    � 9 �A�TD��&$o�3f��T|7�AQxSA`IP����-ø@ T0 k� �S��W�%e1d  3Ab5p�  ��(    � 9 �A�TD��'$o�Cf��T|7�AQxSA`IP����-ü@ T0 k� �S��W�%e1d  3Ab5p�  ��(    � 9 �A�TD��($o�Cf��T|7�AQxSA`IP����-ü@ T0 k� �O��S�%e1d  3Ab5p�  ��(    � 9 �A�TD��($o�Cf��T|7�AQxSA`IP����-ü@ T0 k� �O��S�%e1d  3Ab5p�  ��(   � 9 �A�TD��)$o�Cf��T|7�AQxSA`IP����.ü
@ T0 k� �K��O�%e1d  3Ab5p�  ��(    � 9 �A�TD��+$o�Cf��T|7�AQxSA`IP����.ü
@ T0 k� �K��O�%e1d  3Ab5p�  ��(    � 9 �A�TD��,$o�Cf¸T|7�AQxSA`IP����.ü
@ T0 k� �G��K�%e1d  3Ab5p�  ��(    � 9 �A�TD��-$o�Cf¸T|7�AQxSA`IP����.ü
@ T0 k� �G��K�%e1d  3Ab5p�  ��(    � 9 �A�TD��.$o�Cf¸T|7�AQxSA`IP����.��
@ T0 k� �G��K�%e1d  3Ab5p�  ��(    � 9 �A�TD��/$o�Cf¸T|7�AQxSA`IP����.��
@ T0 k� �G��K�%e1d  3Ab5p�  ��(    � 9 �A�TD��0$o�Cf¸T|7�AQxSA`IP����/��
@ T0 k� �G��K�%e1d  3Ab5p�  ��(    � 9 �A�TD��2$o�Cf¸T|7�AQxSA`IP����/��
@ T0 k� �C��G�%e1d  3Ab5p�  ��(    � 9 �A�TD��3$o�Cf¸T|7�AQxTA`IP����/��	@ T0 k� �C��G�%e1d  3Ab5p�  ��(    � 9 �A�TD��4$o�Cf¸T|7�AQxTA`IP����/��	@ T0 k� �?��C�%e1d  3Ab5p�  ��(    � 9 �A�TD��6$o�Cf¸T|7�AQxTA`IP����/��	@ T0 k� �?��C�%e1d  3Ab5p�  ��(    � 9 �A�TD��7$o�Cf¸T|7�AQtTA`IP����/��	@ T0 k� �?��C�%e1d  3Ab5p�  ��(    � 9 �A�TD��9$o�Cf¸T|7�AQtTA`IP����/��	@ T0 k� �;��?�%e1d  3Ab5p�  ��(    � 9 �A�TD��:$o�Cf¸T|7�AQtTA`IP����0��	@ T0 k� �;��?�%e1d  3Ab5p�  ��(    � 9 �A�TD��;$o�Cf¸T|7�AQtTA`IP����0��	@ T0 k� �7��;�%e1d  3Ab5p�  ��(    � 9 �A�TD��=$o�Cf¸T|7�AQtTA`IP���0��	@ T0 k� �7��;�%e1d  3Ab5p�  ��(    � 9 �A�TE��?$o�Cf¸T|7�AQtTA`IP���0��@ T0 k� �7��;�%e1d  3Ab5p�  ��(    � 9 �A�TE��@$o�Cf¸T|7�AQtTA`IP���0��@ T0 k� �3��7�%e1d  3Ab5p�  ��(    � 9 �A�TE��B$o�Cf¸T|7�AQtTA`IP{���0��@ T0 k� �3��7�%e1d  3Ab5p�  ��(    � 9 �A�TE��C$o�Cf¸T|7�AQtTA`IP{���0��@ T0 k� �3��7�%e1d  3Ab5p�  ��(    � 9 �A�TE��E$o�Cf¸T|7�AQtTA`IP{���1��@ T0 k� �/��3�%e1d  3Ab5p�  ��(    � 9 �A�TF�E$o�Cf¸T|7�AQtTA`IPw���1��@ T0 k� �/��3�%e1d  3Ab5p�  ��(    � 9 �B�*B��� $��s�|7�C�DD�C�D��p�
@ T0 k� �L�P%e1d  3Ab5p�  ��" 	  ��� �B�+B�ǥ $� �{�|7�C�CD�K�D��t�@ T0 k� �P�T%e1d  3Ab5p�  ��" 	  ��� �B� ,B�˥ $�(���|7�C�AD�W����t�@ T0 k� �T�X%e1d  3Ab5p�  ��" 	  ��� �B�(.B�ӥ %�0���|7�C!�@D�_����x�@ T0 k� �\�`%e1d  3Ab5p�  ��" 	  ��� �B�,/B�ۥ %�8���|7�C!�?D�g����|�@ T0 k� �`�d%e1d  3Ab5p�  ��" 	  ��� �B�40B��  %�@���|7�C!�>D�s����| ��@ T0 k� �d�h%e1d  3Ab5p�  ��" 	  ��� �B�81B�� $&�H���|7�C!�=D�{����� ��@ T0 k� �l�p%e1d  3Ab5p�  ��" 	  ��� �B�@2B�� (&�P���|7�C!�;D������ ��@ T0 k� �p �t %e1d  3Ab5p�  ��" 	  ��� �B�D3B��� 0&�T���|7�C!�:D������ ��@ T0 k� �t �x %e1d  3Ab5p�  ��" 	  ��� �B�L4B�� 4'�\���|7�C!�9D������	 ��@ T0 k� �x �| %e1d  3Ab5p�  ��" 	  ��� �B�T5B�� 8'�dϿ�|7�I1�8D�����ΐ
 ��@ T0 k� �|!��!%e1d  3Ab5p�  ��" 	  ��� �B�X6B�� <'�l�Ǽ|7�I1�7D�����Δ
 ��@ T0 k� ��!��!%e1d  3Ab5p�  ��" 	  ��� �B�`7B�� @'�t�ϼ|7�I1�6D�����Θ ��@ T0 k� ��!��!%e1d  3Ab5p�  ��" 	  ��� �B�h8B�'� D(�|�׼|7�I2 5D����Μ ��@ T0 k� ��"��"%e1d  3Ab5p�  �"   ��� B�l9B�/� H(���߼|7�I24D�����Τ ��@ T0 k� Ì"��"%e1d  3Ab5p�  ��/   ��� B�t:B�7�P(����|7�I23D�����Ψ ��@ T0 k� Ð"��"%e1d  3Ab5p�  ��/   ��� B�|;B�C�T)����|7�IB2E���C�ά ��@ T0 k� Ð"��"%e1d  3Ab5p�  ��/   ��� B��<B�K�X)�����|7�IB1E���C�δ ��@ T0 k� Ô"��"%e1d  3Ab5p�  ��/   ��� B��=B�S�\)����|7�IB0E���C��θ ��@ T0 k� Ô"��"%e1d  3Ab5p�  ��/   ��� B��>B�g�h*����|7�IB$/E���C���� �@ T0 k� Ø"��"%e1d  3Ab5p�  ��/   ��� Bќ?B�o�l*͸��|7�I2,.E��C���� �@ T0 k� ��!��!%e1d  3Ab5p� ��/   ��� BѤ@B�w�t*���#�|7�I20.E� C���� �@ T0 k� ��!��!%e1d  3Ab5p� ��/   ��� BѨAB��x*���+�|7�I24-E������ �@ T0 k� ��!��!%e1d  3Ab5p� ��/   ��� BѰBB�|*���3�|7�I28-E������ �@ T0 k� ��!��!%e1d  3Ab5p�  ��/   ��� BѸCB��+���;�|7�I2<,Er ÿ��� �@ T0 k� ��!��!%e1d  3Ab5p�  ��/   ��� E��CB��+���C�|7�IB<,Er(û��� �@ T0 k� ��!��!%e1d  3Ab5p�  ��/   ��� E��DE����+���K�|7�IB@,Er4ó��� �@ T0 k� ��!��!%e1d  3Ab5p�  ��/   ��� E��EE����+���S�|7�IBD+Er<ï��� �@ T0 k� ��!��!%e1d  3Ab5p�  ��/   ��� E��FE���#�,���[�|7�IBH+ErDë�� �@ T0 k� ��!��!%e1d  3Ab5p�  ��/   ��� E��FE���#�,���c�|7�IBH+ErL	ã�� �@ T0 k� ��!��!%e1d  3Ab5p�  ��/   ��� E��GE�Ǧ#�,��k�|7�I2L+ErTß�� �@ T0 k� ��!��!%e1d  3Ab5p�  ��/   ��� E��HE�Ϧ#�,��s�|7�I2P*Er\Û�� �@ T0 k� ��!��!%e1d  3Ab5p�  ��/   ��� E��IE�צ#�,��{�|7�I2P*Er`×��  �@ T0 k� ��!��!%e1d  3Ab5p�  $�/   ��� E��IE��#�-����|7�I2T*Erhӏ��, �@ T0 k� ô"��"%e1d  3Ab5p�  ��/   ��� E��JE��#�-�$���|7�I2T*EbpӋ��4 �@ T0 k� ô"��"%e1d  3Ab5p�  ��/   ��� E�KEr�#�-�,���|7�IBT*EbxӃ��< �@ T0 k� ô#��#%e1d  3Ab5p�  ��/   ��� E�LEs�#�-�8���|7�IBX*Eb��w��L �@ T0 k� ô$��$%e1d  3Ab5p�  ��/   ��� E�MEs��.�@���|7�IBX*Eb��s��T �@ T0 k� ��$��$%e1d  3Ab5p�  ��/   ��� E MEs��.�H���|7�IB\*Eb��k��` �@ T0 k� ��%��%%e1d  3Ab5p�  ��/   ��� E(NEs��.�P���|7�I2\*Eb��g��h �@ T0 k� ��%��%%e1d  3Ab5p�  ��/   ��� E0NEs#��.�X�Ǽ|7�I2\*Eb��_��p �@ T0 k� ��&��&%e1d  3Ab5p�  ��/   ��� E8OEs+��.�`�ϼ|7�I2\*Eb��W��|  �@ T0 k� ��&��&%e1d  3Ab5p�  $�/   ��� E<PEs3��/�h�׼|7�I2\*E��S���  �@ T0 k� 3�'��'%e1d  3Ab5p�  ��/   ��� EDPD�;��/�p�߼|7�I2\*E�!�K���! �@ T0 k� 3�'��'%e1d  3Ab5p�  ��/   ��� E�LQD�C��.�x��|7�IB\*E�"�C���! � @ T0 k� 3�(��(%e1d  3Ab5p�  ��/   �   E�TQD�K��-�|��|7�IB\*E�$�?���" � @ T0 k� 3�(��(%e1d  3Ab5p�  ��/   �   E�\RD�S��,�����|7�IB\*E�&�7���" � @ T0 k� 3�)��)%e1d  3Ab5p�  ��/   �  E�dRD�[��+�����|7�IB\*E�(�/���# �!@ T0 k� ��)��)%e1d  3Ab5p�  ��/   �  E�hREs_��*��	�|7�IB\*E��)�+���# �!@ T0 k� ��*��*%e1d  3Ab5p�  ��/   �  E�pSEsg��)��	�|7�@b\*E��+�#���# �!@ T0 k� ��*��*%e1d  3Ab5p�  ��/   �  E�xSEso�� (��	�|7�@b\*E��-����$ �!@ T0 k� ��+��+%e1d  3Ab5p�  ��/   �  E��SEss��('��	�|7�@b\*E��/����$ �"@ T0 k� ��+��+%e1d  3Ab5p�  $�/   �  E��SEs{��0&��	#�|7�@b\*E��1����% �"@ T0 k� ��,��,%e1d  3Ab5p�  ��/   �  E��SEs���8%��	+�|7�@b\*E��3����% �"@ T0 k� ��-��-%e1d  3Ab5p�  ��/   �  E��TEs���<$��	!/�|7�@b\*E��5�����& �#@ T0 k� ��-��-%e1d  3Ab5p�  ��/   �  E�TEs���D#��	!7�|7�@b\*E��7�����& �#@ T0 k� ��.��.%e1d  3Ab5p�  ��/   �  E�TEc���L#��	!;�|7�@\*E��9����& �#@ T0 k� ��.��.%e1d  3Ab5p�  ��/   �  E�TEc���T"��	!C�|7�@\*E��;����' �#@ T0 k� ��/��/%e1d  3Ab5p�  ��/   �  E�TEc���\!��	!G�|7�@\*Dr�?����' �$@ T0 k� ��0��0%e1d  3Ab5p�  ��/   �  E�TEc���d ��	K�|7�@\*Dr�C���� ( Ӡ$@ T0 k� ��0��0%e1d  3Ab5p�  ��/   �  E�TEc���h��	S�|7�@\*Dr�F����(( Ӡ$@ T0 k� ��1��1%e1d  3Ab5p�  ��/   � 	 E�TEc���p��	W�|7�@\*Dr�H����4( Ӡ$@ T0 k� ��2��2%e1d  3Ab5p�  �/   � 
 S�VEc���x� 	[�|7�@\*Dr�J����<) Ӡ%@ T0 k� ��2��2%e1d  3Ab5p�  ��/   � 
 S�XEc��Ā�	_�|7�@\*Or�L���D) Ӡ%@ T0 k� ��3��3%e1d  3Ab5p�  ��/   �  S�ZEc���|�	!c�|7�@\*Or�N���P* Ӡ%@ T0 k� ��4��4%e1d  3Ab5p�  ��/   �  S�\Ec���|�	!g�|7�@\*Or�P���X* Ӡ%@ T0 k� ��4��4%e1d  3Ab5p�  ��/   �  S�^Ec���x�	!k�|7�@\*OsR���`* Ӝ&@ T0 k� ��5��5%e1d  3Ab5p�  ��/   �  S�`Ec���x�$	!o�|7�@\*OsT���l+ Ӝ&@ T0 k� ��5��5%e1d  3Ab5p�  ��/   �  S�bEc���x�,	!o�|7�@\*OsV	����t+Ӝ&@ T0 k� ��6��6%e1d  3Ab5p�  ��/   �  S�cES���t�4	s�|7�BB\*OsX	����|+Ӝ&@ T0 k� ��7��7%e1d  3Ab5p�  ��/   �  S"�eES���t�<	w�|7�BB\*OsY	���Ј,Ӝ&@ T0 k� ��7��7%e1d  3Ab5p�  ��/   �  S"�gES���t�D	w�|7�BB\*Os[	���А,Ӝ&@ T0 k� ��8��8%e1d  3Ab5p�  ��/   �  S"�hES���p�L	{�|7�BB\*Os ]	���И,Ӡ&@ T0 k� ��9��9%e1d  3Ab5p�  ��/   �  S"�jES���p�T	�|7�BB\*Os$_	��Ф-Ӡ'@ T0 k� ��9��9%e1d  3Ab5p�  ��/   �  S"�lES���p�\��|7�A�\*Os(`	�w�Ь-Ӡ'@ T0 k� ��:��:%e1d  3Ab5p�  ��/   �  S"�mES���p�d���|7�A�\*Os,b	�s���-Ӡ(@ T0 k� ��:��:%e1d  3Ab5p�  ��/   �  S# oES��tp�h���|7�A�\*Os0d	�o���.Ӡ(@ T0 k� ��;��;%e1d  3Ab5p�  ��/   �  S3pES��tp�p���|7�A�\*Os4e	�k���.Ӡ)@ T0 k� ��<��<%e1d  3Ab5p�  ��/   �  S3rES��tp�x���|7�A�\*Os8g	�g���.Ӡ*@ T0 k� ��<��<%e1d  3Ab5p�  ��/   �  S3sES��tl߀���|7�P�\*Os<h	�c���.Ӡ*@ T0 k� ��=��=%e1d  3Ab5p�  ��/   �  S3uEC��tl߈���|7�P�\*Os@j	�_���/Ӡ+@ T0 k� ��>��>%e1d  3Ab5p�   �/   �  S3xEC��tlߘ���|7�P�\*OsHi	�W���/Ӡ-@ T0 k� ��?� ?%e1d  3Ab5p�  ��/   �  S3yEC��tlߠ���|7�P�\*OsLi	�S�� 0Ӡ.@ T0 k� � ?�?%e1d  3Ab5p�  ��/   �  S3{EC��tl
�����|7�P�\*OsPh	�O��0Ӥ/@ T0 k� � @�@%e1d  3Ab5p�  ��/   �  S3|EC��dl	�����|7�P�\*OsTh	�K��0Ӥ1@ T0 k� �A�A%e1d  3Ab5p�  ��/   �  S3 |EC��dl�����|7�P�\*OsXh	�G��0Ӥ2@ T0 k� �A�A%e1d  3Ab5p�  ��/   �  S3${EC��dl�����|7�P�\*F\g	�G��$1Ӥ3@ T0 k� �B�B%e1d  3Ab5p�  ��/   �  S3({E3��dh�����|7�P�\*F`g	�C��01Ӥ5@ T0 k� �B�B%e1d  3Ab5p�  ��/   �  S3,zE3��dh�����|7�P�\*Fhg	�?��D13�8@ T0 k� �D�D%e1d  3Ab5p�  ��/   �  S30zE3��dh �����|7�P�\*Flg	�;��L23�9@ T0 k� �D�D%e1d  3Ab5p�  ��/   �  S34zE3��dk������|7�P�\*Fpg	�;��T23�;@ T0 k� �E�E%e1d  3Ab5p�  ��/   �  S34zCC��dk������|7�P�\*Ftf	�7��`23�<@ T0 k� �F�F%e1d  3Ab5p�  ��/   �  S38yCC��dg������|7�P�\*Fxf	�7��h23�=@ T0 k� �F�F%e1d  3Ab5p�  ��/   �  S3<yCC��dg������|7�P�\*F�g	�3��p3�>@ T0 k� �G�G%e1d  3Ab5p�  ��/   �  S3@yCC��dg�� ���!�7�BB\*E��g	�3��|3�?@ T0 k� �G�G%e1d  3Ab5p�  ��/   �  S3@xCC��Tg�����!�7�BB\*E��g	�3���3�@@ T0 k� �H�H%e1d  3Ab5p�  ��/   �   S3DxCC��Tg�����!�7�BB\*E��g	�3���3�A@ T0 k� �I� I%e1d  3Ab5p�  ��/   � ! S3DxCC��Tg�����!�7�BB\*E��g	�/���3�B@ T0 k� �I� I%e1d  3Ab5p�  ��/   � ! S3HwCC��Tk�� ���!�7�BB\*E��g	�/���4�B@ T0 k� �J� J%e1d  3Ab5p�  ��/   � " S3LwCC��Tk��(���!�7�@\*E��g	�/���4�C@ T0 k� � J�$J%e1d  3Ab5p�  ��/   � " S3LwCS��Tk��0���!�7�@\*E��g	�/���4 �C@ T0 k� � K�$K%e1d  3Ab5p�  ��/   � # S3PwCS��Tk��8���!�7�@\*E��g	�/���4 �C@ T0 k� �$L�(L%e1d  3Ab5p�  ��/   � $ S3TvCS��To��@���!�7�@\*E��g	�/���5 �C@ T0 k� �$L�(L%e1d  3Ab5p�  ��/   � $ S3TvCS��Do��H���!�7�@\*E��g�/���5 �C@ T0 k� �(M�,M%e1d  3Ab5p�  ��/  � % S3XvCS��Do��L���!�7�@\*E��g�/���5 �C@ T0 k� �(M�,M%e1d  3Ab5p�  ��/   � % S3XvCS��Do��T���|7�@b\*E��g�/���5 �C@ T0 k� �,N�0N%e1d  3Ab5p�  ��/   � & S3\uCS��Ds��\���|7�@b\*E��g�/���5 �C@ T0 k� �,N�0N%e1d  3Ab5p�  ��/   � & S3\uCS��Ds��dѿ�|7�@b\*E��g�/���6 �C@ T0 k� �0O�4O%e1d  3Ab5p�  ��/   � ' S3`uCS��Ds��lѿ�|7�@b\*E��g�/���6 �B@ T0 k� �0P�4P%e1d  3Ab5p�  ��/   � ( S3dtCS��Dw��|ѻ�|7�B�`*E�g�/��6 �A@ T0 k� �4Q�8Q%e1d  3Ab5p�  ��/   � ) S3htCc��Dw���ѻ�|7�B�`*E�g�/��6 �A@ T0 k� �4Q�8Q%e1d  3Ab5p�  ��/   � ) S3htCc��Dw���ѷ�|7�B�`*E�f�/��$6 �@@ T0 k� �8R�<R%e1d  3Ab5p�  ��/  � * S3ltCc��4w��ѷ�|7�B�d*E�fB/��,7 �?@ T0 k� �8S�<S%e1d  3Ab5p�  ��/   � + S3ltCc��4{� �	��|7�B�d*EfB/��47 �>@ T0 k� �<S�@S%e1d  3Ab5p�  ��/   � + S3psCc��4{� �	��|7�B�h*IfB/��@7 �=@ T0 k� �<T�@T%e1d  3Ab5p�  ��/   � , S3psCc��4{� �
��!�7�B�h*IfB/��@7 �<@ T0 k� �@T�DT%e1d  3Ab5p�  ��/   � , S3tsCc��4{� �
��!�7�B�l)IfB/��H8 �;@ T0 k� �@U�DU%e1d  3Ab5p�  ��/   � - S3tsCc�� d{� ���!�7�B�p)If�/��P8 �:@ T0 k� �@V�DV%e1d  3Ab5p�  ��/   � . S3xsCc�� d�����!�7�Et)I$f�3��X8 �9@ T0 k� �DV�HV%e1d  3Ab5p�  ��/   � . S3xrCc�� d�����!�7�Ex(I$0f�3��l9 �6@ T0 k� �HW�LW%e1d  3Ab5p�  ��/   � / S3|rCs�� d�����!�7�E|(I$4f�3��t: #�5@ T0 k� �HX�LX%e1d  3Ab5p�  ��/   � 0 S3|rCs�� �������!�7�E�(I$8f�7��|: #�3@ T0 k� �LX�PX%e1d  3Ab5p�  ��/   � 0 S3�rCs�� �������!�7�E�'I$8f�7���: #�2@ T0 k� �LY�PY%e1d  3Ab5p�  ��/   � 1 S3�qCs�� �������!�7�E�'I$8e�;���; #�0@ T0 k� �PZ�TZ%e1d  3Ab5p�  ��/   � 2 S3�qCs�� �������!�7�E�'I8d�;���; #�/@ T0 k� �PZ�TZ%e1d  3Ab5p�  ��/   � 2 S3�qCs�� �������|7�E��&I8d�?���<3�-@ T0 k� �P[�T[%e1d  3Ab5p�  ��/   � 3 S3�qCs��T������|7�E��&I8c�C���<3�,@ T0 k� �T[�X[%e1d  3Ab5p�  ��/  � 3 S3�qCs��T������|7�E��&I8c�G���=3�)@ T0 k� �X\�\\%e1d  3Ab5p�  ��/   � 4 S3�pCs��T�����|7�E��&I$8b�K���=3�(@ T0 k� �`^�d^%e1d  3Ab5p�  ��'   � 5 S3�pCs��T����{�|7�DҰ&I$8b�K���>�&@ T0 k� �h_�l_%e1d  3Ab5p�  ��'   � 6 S3�pCC��T��� �{�|7�DҴ&I$8b�O���>�%@ T0 k� �l_�p_%e1d  3Ab5p�  ��'   � 7 S3�pCC��d���$�w�|7�DҸ&I$8a�S���>�$@ T0 k� �p_�t_%e1d  3Ab5p�  ��'   � 8 S3�pCC��d���,�s�|7�D��&I$8a�W���>�"@ T0 k� �t_�x_%e1d  3Ab5p�  ��'   � 9 S3�pCC��d���0�s�|7�D��&I8a�[�	�?�!@ T0 k� �x_�|_%e1d  3Ab5p�  ��'   � 9 S3�oCC��d���8�o�|7�D��&I8a�_�	�?Ӥ @ T0 k� �x_�|_%e1d  3Ab5p�  ��'   � 9 S3�oCC��d��A<�k�|7�D��'I8a�c�	 ?Ӭ@ T0 k� �x_�|_%e1d  3Ab5p�  ��'   � 9 S3�oCC��d��AD�k�|7�D��'I8a�g�	?Ӱ@ T0 k� �x_�|_%e1d  3Ab5p�  ��'   � 9 S3�oCC��d��AHg�|7�D��'I8a�k�	?Ӵ@ T0 k� �x_�|_%e1d  3Ab5p�  ��'   � 9 S3�oCCǿd��APg�|7�E��'I$8a�o�	#?Ӹ@ T0 k� �x_�|_%e1d  3Ab5p�  ��'   � 9 S3�oCCǽd��ATc�|7�E��(I$8a�w�	#?Ӽ@ T0 k� �x_�|_%e1d  3Ab5p�  ��'   � 9 S3�oE3ǼT��A\!c�|7�E��(I$8a�{�	# ?��@ T0 k� �x_�|_%e1d  3Ab5p�  ��'   � 9 S3�nE3ǺT��A`"_�|7�E��)I$8a��	#(?��@ T0 k� �x_�|_%e1d  3Ab5p�  ��'   � 9 S3�nE3ǶT��Al%�_�|7�E� )@�8a���	4?��@ T0 k� �d[�h[%e1d  3Ab5p�  ��'   � 9 S3�nE3ǵT��Ap&�[�|7�E�*@�8a���	8?��@ T0 k� �TX�XX%e1d  3Ab5p�  ��'   � 9 S3�nE3ǳ���At'�[�|7�E�*@�8a���	<?��@ T0 k� �<U�@U%e1d  3Ab5p�  �'   � 9 �S3�nE3Ǳ���A|)�[�|7�E�+@�8a���	D?��@ T0 k� �$Q�(Q%e1d  3Ab5p�  ��/   � 9 �S3�nE3ǯ���Q�*�[�|7�E�,@�8a���	H?��@ T0 k� �M�M%e1d  3Ab5p�  ��/   � 9 �S3�mE3ǭ���Q�+�[�|7�E� ,G8a���	#L?��@ T0 k� ��J��J%e1d  3Ab5p�  ��/   � 9 �S3�mE3ǫ���Q�-�[�|7�Es(-G8a���	#P?��@ T0 k� ��F��F%e1d  3Ab5p�  ��/   � 9 �S3�mE3ǧė�Q�0�[�|7�Es4/G8a���	#X?��@ T0 k� ��?��?%e1d  3Ab5p�  �/   � 9 �S3�mISǥė�Q�1�_�|7�Es</G8a���	#\?��@ T0 k� ð?��?%e1d  3Ab5p�  ��/   � 9 �S3�mISǣė�	Q�3�_�|7�Es@0G8a���	`?��@ T0 k� ô@��@%e1d  3Ab5p�  ��/   � 9 �S3�mISǡē�	Q�4�_�|7�Es@0G8a���	d?��@ T0 k� ô@��@%e1d  3Ab5p� ��/   � 9 �S3�mISǠē�	Q�5�_�|7�I�D1G8a���	h@��@ T0 k� ø@��@%e1d  3Ab5p� ��/   � 9 �S3�lISǜԓ�	Q�8�c�|7�I�L1G8a���	p@��@ T0 k� ��A��A%e1d  3Ab5p� ��/   � 9 �S3�lIcǛԓ�	Q�9�c�|7�I�P1G$8a���	#tA3�@ T0 k� ��B��B%e1d  3Ab5p� ��/   � 9 �S3�lIcǙԏ�	a�:�g�|7�I�X2G$8a���	#xA3�@ T0 k� ��B��B%e1d  3Ab5p� ��/   � 9 �S3�lIcǘԏ�	a�;�g�|7�I�\2G$8a���	#|A3�@ T0 k� ��B��B%e1d  3Ab5p� ��/   � 9 �S3�lIcǖԋ�	a�<�g�|7�I�\2G$8a���	#�A3�@ T0 k� ��C��C%e1d  3Ab5p� ��/   � 9 �S3�lIcǕԋ�	a�=�k�|7�I�`2G$8a���	#�A3�@ T0 k� ��C��C%e1d  3Ab5p� ��/   � 9 �S3�lISǔԇ�	a�>�k�|7�I�d2G$8a���	�B3�@ T0 k� ��D��D%e1d  3Ab5p� ��/   � 9 �S3�lISǒ��	Q�>�o�|7�I�h2G$8a��	�B3�@ T0 k� ��D��D%e1d  3Ab5p� ��/   � 9 �S3�lISǑ��	Q�?�s�|7�I�l2G$8a��	�B3�@ T0 k� ��C��C%e1d  3Ab5p� ��)   � 9 �S3�kISǏ�{�	Q�A�w�|7�E�p3G$8a��	�B3�@ T0 k� ��B��B%e1d  3Ab5p� ��)   � 9 �S3�kIcǎ�{�	Q�B�w�|7�E�t3G$8a��	#�B3�@ T0 k� ��A��A%e1d  3Ab5p� ��)   � 9 �S3�kIcǍ4w�!�C�{�|7�E�x3G$8a��	#�B��@ T0 k� ��A��A%e1d  3Ab5p� ��)   � 9 �S3�kIcǌ4s�!�D�|7�E�x3G$8a�  	#�B��@ T0 k� ��A��A%e1d  3Ab5p� ��)   � 9 �S3�kIcǋ4s�!�E�|7�E�x3G$8a�$	#�B��@ T0 k� ��A��A%e1d  3Ab5p� ��)   � 9 �S3�kIcǉ4o�!�G��|7�Ec|3G$8a�,	#�B��@ T0 k� ��A��A%e1d  3Ab5p� ��)   � 9 �SC�kISÊTo�!�H��|7�Ec�3G$8a�0	�C��@ T0 k� �A��A%e1d  3Ab5p� ��)   � 9 �SC�kISÊTo�!�I��|7�Ec�3G$8a�4	�C��@ T0 k� �A��A%e1d  3Ab5p� ��)   � 9 �SC�kISÊTo��J��|7�Ec�4G$8a�8	�C��@ T0 k� �A��A%e1d  3Ab5p� ��)   � 9 �SC�kISÊTo��K��|7�Ec�4G$8a�<	�C��@ T0 k� �A��A%e1d  3Ab5p� ��)   � 9 �SC�jISÊTo��L��|7�Ec�4G$8a�@		�C��@ T0 k� �A��A%e1d  3Ab5p� ��)   � 9 �SC�jASÊTs��M��|7�ES�4G$8a�D
	#�C��@ T0 k� ��A��A%e1d  3Ab5p� ��)   � 9 �SC�jASËTs��O��|7�ES�4@�8a�D	#�C��@ T0 k� ��A��A%e1d  3Ab5p� ��)   � 9 �SC�jASËTs� P��|7�ES�4@�8a�H	#�C��@ T0 k� ��A��A%e1d  3Ab5p� ��)   � 9 �SC�jAS��Ts�Q��|7�ES�4@�8a�L	#�C��@ T0 k� ��A��A%e1d  3Ab5p� ��)   � 9 �U�jAS��Tw�R��|7�ES�4@�8a�L	#�C��@ T0 k� ��A��A%e1d  3Ab5p�  ��)   � 9 �U�jE㿋Tw�S��|7�A�5@�8a�P	�C��@ T0 k� �A��A%e1d  3Ab5p�  ��)   � 9 �U�jE㻋Tw�S��|7�A�5@d8a�P	�C��@ T0 k� �A��A%e1d  3Ab5p�  .�)   � 9 �U�jE㻌Tw�T��|7�A�5@d8a�T	�C��@ T0 k� �A��A%e1d  3Ab5p�  ��)   � 9 �U�jE㷌Tw��U��|7�A�5@d8a�T	�C��@ T0 k� �A��A%e1d  3Ab5p�  ��)   � 9 �U�jE㷌T{��$V��|7�A�5@d8a�T	�C��@ T0 k� �A��A%e1d  3Ab5p�  ��)   � 9 �U�jE�T{��(W��|7�A|4@d8a�T�C��@ T0 k� ��E��E%e1d  3Ab5p�  ��)   � 9 �U�jE�T{��0X��|7�A|4@8a�T�C��@ T0 k� ��A��A%e1d  3Ab5p�  �)   � 9 �U�jE�T{��4X��|7�C�|4@8a�X�C��@ T0 k� ��<��<%e1d  3Ab5p�  ��/   � 9 �@c�iE�T{��<Y��|7�C�x4@8a�X�C��@ T0 k� ��8��8%e1d  3Ab5p�  ��/   � 9 �@c�iE�T{��@Z��|7�C�x4@8a�X�C��@ T0 k� ��3��3%e1d  3Ab5p�  ��/   � 9 �@c�iE�T��HZ���|7�C�t4@8a�Xc�C��@ T0 k� ��/��/%e1d  3Ab5p�  ��/   � 9 �@c�iF��T��L[���|7�C�t3@�8a�Tc�C��@ T0 k� �p*�t*%e1d  3Ab5p�  �/   � 9 �@c�iF��T��T[���|7�E�p3@�8aSTc�C�@ T0 k� �p*�t*%e1d  3Ab5p�  ��/   � 9 �E��hF��T��X[���|7�E�p3@�8aSTc�C�@ T0 k� �t*�x*%e1d  3Ab5p� ��/   � 9 �E��hF��T�r`\���|7�E�l3@�8aST c�C�@ T0 k� �t*�x*%e1d  3Ab5p� ��/   � 9 �E��gF��T�rl\	�|7�E�d3@�8aSP"s�C�@ T0 k� �x)�|)%e1d  3Ab5p� ��/   � 9 �E��gF��T�rp\	�|7�E�d3@�8aCP#s�C�@ T0 k� �x)�|)%e1d  3Ab5p� ��/   � 9 �E��fF��T��rx\	�|7�E�d3A8aCL#s�C�@ T0 k� �|)��)%e1d  3Ab5p� ��/   � 9 �E��fF��T��r|\	�|7�C�`4A8aCL#s�C�@ T0 k� �|)��)%e1d  3Ab5p� ��/   � 9 �E��eF��T��r�\	�|7�C�\4A8aCL$s�C�@ T0 k� Ӏ(��(%e1d  3Ab5p� ��/   � 9 �E��eF��T��r�\	"�|7�C�X5A8aCH$��C�@ T0 k� Ӏ(��(%e1d  3Ab5p� ��/   � 9 �E��dF��T��r�\	"�|7�C�T5A8aCH$��C�@ T0 k� ӄ(��(%e1d  3Ab5p� ��/   � 9 �E��dF��T��r�\	"�|7�C�T6AT8aCH$��C�@ T0 k� �(��(%e1d  3Ab5p� ��/   � 9 �E��cF��T��r�\	"#�|7�C�P6AT8aCD%��C�@ T0 k� �'��'%e1d  3Ab5p�  ��/   � 9 �E��bF��T��r�\	"#�|7�C�L7AT8aCD%��C�@ T0 k� �'��'%e1d  3Ab5p�  ��/   � 9 �E��aF��T��b�[	'�|7�C�D7AT8aCD%��C�@ T0 k� �'��'%e1d  3Ab5p�  ��/   � 9 �E��aF��T��b�[	+�|7�C�@8AT8aCD%��C�@ T0 k� �'��'%e1d  3Ab5p�  ��/   � 9 �E��`F��T��b�Z	+�|7�C�<8C�4aCD%��C�@ T0 k� �'��'%e1d  3Ab5p�  ��/   � 9 �E��_F��T��b�Z	/�|7�C�88C�4aCD%��C�@ T0 k� �&��&%e1d  3Ab5p�  /�/   � 9 �E��^F��T��b�Z	/�|7�C�49C�4aCD%��C�@ T0 k� �&��&%e1d  3Ab5p�  ��/   � 9 �E��]F��T��b�Y	"3�|7�C�09C�0aCD%��C�@ T0 k� �&��&%e1d  3Ab5p�  ��/   � 9 �E��]F��T��b�Y	"3�|7�C�(:C�0aCD%��C�@ T0 k� �&��&%e1d  3Ab5p�  ��/   � 9 �E��\F��T��b�X	"3�|7�C�$:ED,`CD%��C�@ T0 k� �%��%%e1d  3Ab5p�  ��/   � 9 �E��[BC��T��b�W	"7�|7�C�:ED,`CD%��C�@ T0 k� �%��%%e1d  3Ab5p�  ��/   � 9 �E��ZBC��T��R�W	"7�|7�C�;ED(`�D%��C�@ T0 k� �%��%%e1d  3Ab5p�  ��/   � 9 �E��YBC��T��R�V	7�|7�C�;ED$`�D%��C�@ T0 k� �%��%%e1d  3Ab5p�  ��/   � 9 �E��XBC��T��R�V	7�|7�C�;ED$`�D%��C�@ T0 k� �$��$%e1d  3Ab5p�  ��/   � 9 �E��WBC��T��R�U	;�|7�C�<ED _�D%��C�@ T0 k� �$��$%e1d  3Ab5p�  ��/   � 9 �E��VBC��T��R�U	;�|7�C� <ED_�D%�C�@ T0 k� �$��$%e1d  3Ab5p�  ��/   � 9 �E��VA�T��R�T	;�|7�C��=ED_�D%�C�@ T0 k� �$��$%e1d  3Ab5p�  �/    � 9 �C��UA�T��R�T b;�|7�AR�=ED^�D%�C�@ T0 k� �$��$%e1d  3Ab5p�  �/    � 9 �C��TA�T��R�S b;�|7�AR�=A^�D%�C�@ T0 k� �#��#%e1d  3Ab5p�  ��/    � 9 �C��SA�T��R�S b;�|7�AR�>A^�D%�C�@ T0 k� �#��#%e1d  3Ab5p�  ��/    � 9 �C��SA�T��R�R b;�|7�AR�>A]�D$S�C�@ T0 k� �#��#%e1d  3Ab5p�  ��/    � 9 �C��RD���T��R�R b;�|7�AR�>A]�D$S�C�@ T0 k� �#��#%e1d  3Ab5p�  ��/    � 9 �C��QD���T��B�Q �;�|7�AR�?A]�D$S�C�@ T0 k� �"��"%e1d  3Ab5p�  ��/    � 9 �C��QD���T��B�Q �;�|7�AR�?A\�D$S�C�@ T0 k� �"��"%e1d  3Ab5p�  ��/    � 9 �C��QD���T��B�P �;�|7�AR�?A\�D$S�C�@ T0 k� �"��"%e1d  3Ab5p�  ��/    � 9 �C��QD���T��B�P �;�|7�AR�?A \�D$3�B�@ T0 k� �"��"%e1d  3Ab5p�  ��/    � 9 �C��PD���T��B�P �;�|7�AR�@A�[�D$3�B�@ T0 k� �"��"%e1d  3Ab5p�  ��/    � 9 �C�PD���T�� ��PB;�|7�AR�@A�[�D$3�A�@ T0 k� �!��!%e1d  3Ab5p�  ��/    � 9 �C�PD���T�� ��OB;�|7�AR�@A�[�D$3�@�@ T0 k� �!��!%e1d  3Ab5p�  ��/    � 9 �C�PD���T�� ��OB;�|7�AR�AA�Z�D$3�@�@ T0 k� �!��!%e1d  3Ab5p�  ��/    � 9 �C�OD���T�� ��OB?�|7�AR�AA�Z�D$3�?�@ T0 k� �!��!%e1d  3Ab5p�  ��/    � 9 �C�OD���T�� ��OB?�|7�AR�AA�Z�D$3�>�@ T0 k� �!��!%e1d  3Ab5p�  ��/    � 9 �C�OD���T�� ��O"?�|7�AR�AA�Z�D$3�>�@ T0 k� � �� %e1d  3Ab5p�  ��/    � 9 �C�OD���T�� b�O"?�|7�AR�BA�Y�D$3�=�@ T0 k� � �� %e1d  3Ab5p�  ��/    � 9 �C�ND���T�� b�O"?�|7�AR�BA�Y�D$3�<�@ T0 k� �� �� %e1d  3Ab5p�  ��/    � 9 �C�ND���T�� b�O"C�|7�AR�BA�Y�D$C�;�@ T0 k� �� �� %e1d  3Ab5p�  ��/    � 9 �C�ND���T�� b�O"C�|7�AR�CA�X�D$C�:�@ T0 k� ����%e1d  3Ab5p�  ��/    � 9 �C�ND���T�� b�P"C�|7�AR�CA�X�D$C�9�@ T0 k� ����%e1d  3Ab5p�  ��/    � 9 �C�MD���T����P"G�|7�AR�CA�X�D$C|9�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �C�MD���T����P�G�|7�AR�CA�X�D$Cx8s�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �D�MD���T����P�K�|7�AR|DA�W�D$�t7s�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �D�MD���T����P�K�|7�ARxDA�W�D$�t6s�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �D�MD���T����Q�O�|7�ARtDA�W�D$�p5s�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �D|LD���T����Q�O�|7�ARpDA�W�D$�l4s�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �DxLD���T����Q�O�|7�ARhDA�V�D$�h3��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�tLD���T����Q�S�|7�ARdEA�V�D$�d2��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�lLD���T���Q�S�|7�AR`EA�V�D#�d2��@ T0 k� ����%e1d  3Ab5p�  ��*   � 9 �E�hLD���T���Q�W�|7�AR`EA�V�D#�d2��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�dKD���T���Q�W�|7�AR\EA�V�D#�d2��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�\KD���T���Q�X |7�ARXFA�U�D#�d2��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�XKD���T���Q�X|7�ARTFA�U�@"�d2 3�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�PKD���T�� b�QBX|7�ARPFA�U�@"�`1 3�@ T0 k� ��
��
%e1d  3Ab5p�  ��*    � 9 �E�LKD���T�� b�QB\|7�ARLFA�U�@!�`1 3�@ T0 k� ��
��
%e1d  3Ab5p�  ��*    � 9 �E�DKD���T�� b�QB\|7�ARHFA�T�@!�\1 3�@ T0 k� ��
��
%e1d  3Ab5p�  ��*   � 9 �E�@KD���T�� b�QB`|7�ARDGA�T�@ �\0 3�@ T0 k� ��
��
%e1d  3Ab5p�  ��*    � 9 �E�8KD���T�� b�QB`|7�AR@GA�T�< �X0��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�4KD���T����Q"d	|7�AR<GA�T�< �X0��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�,KD���T����Q"d
|7�AR<GA�T�<�X/��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�(KD���T����R"h|7�AR8GA�T�<�T/��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E� KD���T����R"h|7�AR4HA�S�<�T/��@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�LD���T����R"l|7�AR0HA�S�<�T/C�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�LD���T����R"p|7�AR,HA�S�8�P.C�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�LD���T����S"p|7�AR,HA�S�8�P.C�@ T0 k� ����%e1d  3Ab5p�  ��*    � 9 �E�LD���T����T�t|7�AR(HA�S�8�L.C�@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �E�LD���T����U�x|7�AR$HA�R�8�L.C�@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �E�LD���T��"�U�x|7�AR IA�R�8�L-S�@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �E�LD���T��"�V�||7�AR IA�R�8�H-S�@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �D�LEc��T��"�W�|7�ARIA�R�4�H-S�@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �D�LEc��T��"�X��|7�ARIA�R�4�H-S�@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �D� LEc��T��"�Y��|7�ARIA�R�4�D,S�@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �D� LEc��T����Y��|7�ARIA�Q�4�D,S�@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �D��LEc��T����Z��|7�ARJA�Q�4�D,S�@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �D��LEc��T����[��|7�ARJA�Q�4�@,��@ T0 k� ���%e1d  3Ab5p�  ��*   � 9 �D��LEc��T����\��!|7�ARJA�Q�0�@+��@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �D��LEc��T����]��#|7�ARJA�Q�0�@+��@ T0 k� ���%e1d  3Ab5p�  ��*    � 9 �D��LD3��T����]B�$|7�ARJA�Q�0�@+��@ T0 k� �x�|%e1d  3Ab5p�  ��*    � 9 �D��LD3��T����^B�&|7�ARJA�Q�0�<+��@ T0 k� �p�t%e1d  3Ab5p�  ��*    � 9 �D��LD3��T����_B�(|7�AR JA�P�0�<*��@ T0 k� �p�t%e1d  3Ab5p�  ��*    � 9 �D��MD3��T����_B�*|7�AR KA�P�0�<*��@ T0 k� �p�t%e1d  3Ab5p�  ��*    � 9 �D��MD3��T����`B�+|7�AQ�KA�P�0�8*��@ T0 k� �l�p%e1d  3Ab5p�  ��*    � 9 �A��MD3��T����a"�-|7�AQ�KA�P�,�8*��@ T0 k� �h�l%e1d  3Ab5p�  ��*    � 9 �A��MD3��T����b"�/|7�AQ�KA�P�,�8*��@ T0 k� �d�h%e1d  3Ab5p�  ��*    � 9 �A��MD3��T����b"�1|7�AQ�KA�P�,�8)��@ T0 k� �`�d%e1d  3Ab5p�  ��*    � 9 �A��ND3��T��¼c"�3|7�AQ�KA�P�,�4)��@ T0 k� �X�\%e1d  3Ab5p�  �*    � 9 �A��NL3��T��¼d"�4|7�AQ�KA�P�,�4)s�@ T0 k� �L�P%e1d  3Ab5p�  ��/    � 9 �F�NL3��T��¼d"�6|7�AQ�KA�O�,�4)s�@ T0 k� �8�<%e1d  3Ab5p�  ��(    � 9 �F�OL3�T��¼e"�8|7�AQ�LA�O�,�4)s�@ T0 k� �,�0%e1d  3Ab5p�  ��(    � 9 �F�OL3�T��¼e�:|7�AQ�LA�O�(�0(s�@ T0 k� �$�(%e1d  3Ab5p�  ��(    � 9 �F�PL3{�T��¸f�<|7�AQ�LA�O�(�0(s|@ T0 k� �� %e1d  3Ab5p�  ��(    � 9 �F�PL3{�T��¸g��=|7�AQ�LA�O�(�0(sx@ T0 k� ��%e1d  3Ab5p�  ��(    � 9 �F�QL3w�T��¸g��?|7�AQ�LA�Oc(�0(st@ T0 k� �
�
%e1d  3Ab5p�  ��(    � 9 �F�QL3w�T�¸h��A|7�AQ�LA�Oc$�,(�p@ T0 k� ��%e1d  3Ab5p�  ��(    � 9 �F�QL3pT�¸h	2�B|7�AQ�LA�Oc$�,(�l@ T0 k� � �%e1d  3Ab5p�  ��(    � 9 �F�RL3lT�´i	2�D|7�AQ�LA�Oc �,'�h@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�RL3lT�´j	2�E|7�AQ�LA�Nc �,'�h@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�RL3hT�´j	2�E|7�AQ�MA�NS�,'�d@ T0 k� ��	��	%e1d  3Ab5p�  ��(    � 9 �F�RL3hT�´k	2�E|7�AQ�MA�NS�('�`@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�SL3d	T�´k��F!�7�AQ�MA�NS�('�`@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�SLCd�´l��G!�7�AQ�MA�NS�('�`@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�TLC`�°l��H!�7�AQ�MA�NS�$'�`@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�TLC`�°m��H!�7�AQ�MA�Nc�$'s`@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�ULC\�°m��I!�7�AQ�MA�Nc� 's\@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�ULC\�°n��I!�7�AQ�MA�Nc� 's\ @ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�ULC\�°n��J!�7�AQ�MA�Nc�'sX!@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �F�VLCX{�°o��K!�7�AQ�MA�Nc �'sX!@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�VLCX{�°o��K!�7�AQ�NA�Mb��'sX!@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�VLCT{�¬p��K!�7�AQ�NA�Mb��'sX!@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�VLCT{�¬p��K!�7�AQ�NA�Mb��'sX"@ T0 k� ���%e1d  3Ab5p�  ��(   � 9 �F�WLCP{�¬q��K|7�AQ�NA�Mr��'sX#@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�WLCP{�¬q��L|7�AQ�NA�Mr��'sT#@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�WLCP{�¬q��L|7�AQ�NA�Mr��'sT$@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�WLCL{�¬r��L|7�AQ�NA�Mr��'sT%@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�WLCL${�¬r��L|7�AQ�NA�Mr��'sT%@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�WLCH${�¬s��L|7�AQ�NA�Mr��'sP&@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�WLCH${�¨s��M|7�AQ�NA�Mr��'sP&@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �F�WLCH${�¨s��M|7�AQ�NA�Mr��'sP'@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �BB�WLCD${�¨t��M|7�AQ�OA�Mr��(sL(@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �BB�WLCD${�¨t��M|7�AQ�OA�Mr�
�(3L(@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �BB�WLCD${�¨u��M|7�AQ�OA�Lr�
� (3L)@ T0 k� �x�|%e1d  3Ab5p�  ��(    � 9 �BB�WLC@${�¨u��M!�7�AQ�OA|L��
� (3L*@ T0 k� �p�t%e1d  3Ab5p�  ��(    � 9 �BB�WLC@$w�¨u��M!�7�AQ�OA|L��
��(3H*@ T0 k� �d�h%e1d  3Ab5p�  ��(    � 9 �BB�WLC@$w�¨v��N!�7�AQ�OA|L��	��(3H+@ T0 k� �\�`%e1d  3Ab5p�  ��(    � 9 �BB�WLC<$w�¨v��N!�7�AQ�OA|L��	��(�H+@ T0 k� �T
�X
%e1d  3Ab5p�  ��(    � 9 �BB�WLC<$w�¤w��N!�7�AQ�OA|L��	��(�H+@ T0 k� �P
�T
%e1d  3Ab5p�  ��(    � 9 �BB�WLC<$w���w��N!�7�AQ�OA|L����(�D,@ T0 k� �H
�L
%e1d  3Ab5p�  ��(    � 9 �A��WLC8$w���w��O!�7�AQ�OA|L����(�D,@ T0 k� �D
�H
%e1d  3Ab5p�  ��(    � 9 �A��WLC8$w���x��O!�7�AQ�OAxL����(�D,@ T0 k� �<	�@	%e1d  3Ab5p�  ��(    � 9 �A��WLC8$w���x��O!�7�AQ�OAxL����(�D,@ T0 k� �4	�8	%e1d  3Ab5p�  ��(    � 9 �A��WLC4$w���x��O!�7�AQ�OAxL����(�@,@ T0 k� �,	�0	%e1d  3Ab5p�  ��(    � 9 �A��WLC4$w���y��O!�7�AQ�OAxL�x��(�@,@ T0 k� �(	�,	%e1d  3Ab5p�  ��(    � 9 �LR�WLC4$w�"�y��O|7�AQ�PAxL�p��(�@,@ T0 k� � �$%e1d  3Ab5p�  ��(    � 9 �LR�WLC0$w�"�y��O|7�AQ�PAxL�l��(�@,@ T0 k� ��%e1d  3Ab5p�  ��(    � 9 �LR�WLC0$w�"�z��O|7�AQ�PAxL�d��(�@,@ T0 k� ��%e1d  3Ab5p�  ��(    � 9 �LR�WLC0$w�"�y��O|7�AQ�PAxL�\��( C<,@ T0 k� ��%e1d  3Ab5p�  ��(    � 9 �LR�WLC,$w�"�y��P|7�AQ�PAtL�T��( C<,@ T0 k� ��%e1d  3Ab5p�  ��(    � 9 �LR�WLC,$w��y��P|7�AQ�PAtK�L��( C<,@ T0 k� ��� %e1d  3Ab5p�  ��(    � 9 �LR�WLC,$w��y��P|7�AQ�PAtK�D��( C@,@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �LR�WLC($w��x��P|7�AQ�PAtK�<��( C@,@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �LR�WLC($w��x��P|7�AQ�PAtK�8��( C@,@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �LR�WL3($w��x��Q|7�AQ�PAtK�0��( C@+@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �Lb�WL3$$w��x��Q|7�AQ�PAtK�(��( CD+@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �Lb�WL3$$w��w¼Q|7�AQ�PAtKb ��( CD+@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �Lb�WL3$$w��w¼Q|7�AQ�PAtKb��) CD*@ T0 k� ����%e1d  3Ab5p�  ��(    � 9 �Lb�WL3 $w���w¼Q|7�AQ�PAtKb��) CH)@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WL3 $s���w¼R|7�AQ�PApKb��) SL)@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WD3 $s���v¼R|7�AQ�PApKb ��) SL(@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WD3$s���v¼R|7�AQ�PApKQ���) SP(@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WD3$s���v¼R|7�AQ�QApKQ���) SP'@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WD3$s���u¼R|7�AQ�QApKQ���) ST&@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WD3$s���u¼R|7�AQ�QApKQ���)�T&@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WL3$s���t¼S|7�AQ�QApKQ���)�X%@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WL3$s���t��S|7�AQ�QApKQ���)�X%@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WL3$s���s��S|7�AQ�QApKQ���)�\$@ T0 k� ���%e1d  3Ab5p�  ��(    � 9 �Lb�WL3s���r��S|7�AQ�QApKQ���)�\$@ T0 k� �|��%e1d  3Ab5p�  ��(    � 9 �Lb�WL3s���r��S|7�AQ�QApKQ���)�`#@ T0 k� �x�|%e1d  3Ab5p�  ��(    � 9 �Lb�WL3s���q��S|7�AQ�QAlKQ���)�`"@ T0 k� �t�x%e1d  3Ab5p�  ��(    � 9 �Lb�WL3s�r�q��S|7�AQ�QAlKQ���)�d"@ T0 k� �l�p%e1d  3Ab5p�  ��(    � 9 �Lb�WL3s�r�p��T|7�AQ�QAlKQ���)�d!@ T0 k� �h�l%e1d  3Ab5p�  ��(    � 9 �Lb�WL3s�r�o��T|7�AQ�QAlKQ���)�h!@ T0 k� �`�d%e1d  3Ab5p�  ��(    � 9 �Lb�WL3Ts�r�n��T|7�AQ�QAlKQ���)�h @ T0 k� �\�`%e1d  3Ab5p�  ��(    � 9 �Lb�WL3Ts�r�m��T|7�AQ�QAlJQ���)�l @ T0 k� �T�X%e1d  3Ab5p�  ��(    � 9 �Lb�WLCTs���l��T|7�AQ�QAlJQ���)�l@ T0 k� �P�T%e1d  3Ab5p�  ��(    � 9 �Lb�WLCTs���k��T|7�AQ�QAlJQ���)�p@ T0 k� �D �H %e1d  3Ab5p�  ��(    � 9 �Lb�WLCTs���j��T|7�AQ�QAlJQ���)�p@ T0 k� �< �@ %e1d  3Ab5p�  ��(    � 9 �Lb�WLCTs���i��T|7�AQ�QAlJQ���)�t@ T0 k� �8 �< %e1d  3Ab5p�  ��(    � 9 �                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��"t ]�*O*N  �� T��    	  � �9,     T�� �9,    	�   	           	 Z �          �     ���   0
%            EO?  ` `       � ��t     E�X ���    ���   	        ) Z �         ���  �  ���  8	          ��d   � �
	   �q    ��.�q    ��     	          Z �         �`�    ���   0	           f�:   � �	     ��     f�: ��           	           	 Z �          ���    ���   8          T(�   � �
	   . �Ǖ     T(� �Ǖ                     J 	 Z �          � �    ���   P
		         ��z�  ��	     B���    ��z����                             ���l              q  ���    P              T5�        V ]�7     T2O ]��     6��             P��          �`  �  ��@   0           I��       j �P�     I�� �S�      ��               ��          �      ��@   0	
          ��A         ~ �X    �� H    ���            �   �         ��     ��J   0          1+-    	     � ���     1
� ��    ��+            	     �         	 F   �  ��B   0
	          c� ��
      � �'�     ~	 ��    �q�                      �� �       
       E  ��@    		 5            ��H       �  �q    ��H  �q               ��        � !          �@       ��F   8'                 ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��d%  ��        � n�    ��j� þ    ��� "                x                j  �       �                         ��    ��        �       ��              "                                                �                          � � � �� ] �  � �  ��   
 	               
  @    �� �b�A       K� �^@ L�  _@ K�  _� �$  g  �d g@ �� g`���J ����X ����� � ˤ ]` �� ]����. ����< ����J ����X � �� �r` �� s` �� o� �� �o� �� p� 
�| W� 
�\ W� �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �D �Q` � }`���� ����� � 
�| V� 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� �  9���>  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"     
�j,� B �
� �  �  
� ����  ��     �       ����  ��     �      ����  ��     �           � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �(      �� � �  ���        � �T ��        �        ��        �        ��        �  
  ��    ������n        ��                         ��  0 �� ��                                    �                 ����            ��  ���%��   9 ���               �HFD y Yake ne   y   0:00                                                                        3  2     �C
� �@kV` k^ �c� � c� � �C. � C6  C7! �	C8! � 
C: � C; �J� �J� �J� �J� �J� �C' � C"- �C#  �C%( � C'0 �kj �kr � �c� � �c� � � c� � �	� � �	� � �� � �� � xC � x  C � y !C � q "C � i #C � a $C � �%"� � � &"� � �'"� � �(*� � z )*OW z**(_ �+**o �,*8g � -*Gg � .*Ew � /*Pg �0" �1*o 2*Fg3)�w*4*8g: 5*Gg:  *Ew: 7*Gg:  *Ew: 9*JwJ )�g �;)�g �<**=*<g
>*2w* *:g                                                                                                                                                                                                                         �� R         �    @ 
         �     ^ P E a  ������              	 �������������������������������������� ���������	�
��������                                                                                          ��    �`�� ��������������������������������������������������������   �4, 5� * ۂ�@~��@���4�� �������                                                                                                                                                                                                                                                                                                                               @=@���ژ                                                                                                                                                                                                                                             +    ��  D�J    	  �  	                           ������������������������������������������������������                                                                                                                                     |     �      �        �          �     �    	  
 	 
 	 	 ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� �������            �                p    $         K
�J                                     ������������������������������������������������������                                                                                                                                        �      �              ��      ��   �          	 	 
  	 
 
 ��  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���            x                                                                                                                                                                                                                                                                                                   
        �             


             �  }�                                    +!                              '     'u               ����������������   	����������������������������      O������������  +  +����������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" R > / 	              	                  � !ϛ^ �\        �c�b7.P�1sc$                                                                                                                                                                                                                                                               )n)n1n  
�              b            a                  `      m                                                                                                                                                                                                                                                                                                                                                                                                        > �  >�  J�  @�  2�  EZm_  �N U���_��������� ~�˖�l��������������̕        6  ���B : ���         	 	 �   & AG� �  �   
           	A\�                                                                                                                                                                                                                                                                                                                                       B F   h                      !��                                                                                                                                                                                                                            Y��   �� �� ��      �� B 	     ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� ���������  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���      �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    :      :     ��                       B     �  �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��[�  �    � �$ ^$    ����  �}  ޢ  ��  �1   �    >     �f ��        p���� ��   p���� �$     � ���h  �   � ��� �    � �N ^$�V   �  ��"       &����     &h��m ���>�������J s y 
n� ����� ��� �����   � ��� ��  � ��� ` �s �s��   �      �  ��   ����� e�����  g���          f ^�   �      ��� 9      �      ��"����2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "! ""! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                        "!  " ! " ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                      �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �             ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                                                                                                                                                                    �� ������}����zvw� w
�  �� 	�� �� �� ��� �̽ ��� ɪ  ̘ ��,̾�-�� ��                  ��       �                                 ��  ��  ��� ��� �������̼���������˸�˸�+���"��U�X�U�EU�UDH�UTX�U3U�T3E�@3��	��  �� ��"�"""�"""���  ��            �   �   P   T   U   T   S   C   3   30  30  ;�  ��  ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    � ��  �   ��  �                                       "  "  "                                                                                                                                                                      �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��                     ��  ��  ���     �     �                                                                                                                                                                                      �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                �  �  �   �   ��  �                            �   ���                            �   �                                                                                                  "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��  �       �                        �   ��  ���  � �    �                                                                                                                                             �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �          �  � � �� ��     � ��  ��  ɀ  �   ��  ��  ���   �   �   �                                                                                                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                        �          �   � � �  ��� ��  �                       �   �                      �������  ���    �              �  �� ��  �    � ���                                                                                                                                                                                                           �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �   �           �   �             
�  ��  ��  ��  �����  �   �          ��                           � ��                    ���� �                             � �������������  �                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    �   �                             �  ��  ��  ww  ��  vv  w"   "   "  �� ��                   ����������             ��  �   ��  �                             �  �˰ ��� �wp ���                                                                                                                                                                 �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                  �    �                    ��                      �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                    �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  ���" �!  �  �� �   �                  �   �  �  �   �               �   �                     �                        �         �  �� �  �� ��                                                                                                                                       ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r`    /   �  �   ��                             �                        ���� ��� ����                � ��                    ���� �                                                                                                                                                                                                    �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""���������������������""""������II������""""������IIII""""������DI�I�""""������DI�I�""""�����IIDIIIA""""��������DD""""������IADD�A��""""��������I���I�������I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=""""��������AA�A    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ADA�LL��L�D����3333DDDD x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(XxLL����������D����3333DDDD w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""����������A������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(""""�������I�I������ �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�""""�������I��D���I�������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7�D�M�D���M������3333DDDD  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`D�M�A�����MD�����3333DDDD 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
""""�����AMAD������ w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw""""������������������ w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xwwfFfFDfFFfFffdFffff3333DDDD + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+DDFFDfFFfdFffff3333DDDD � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(�""""wwwwwwwGGD � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(�""""wwwwwwqwAqwAwA �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(�""""wwwwqwqAwAqAqAq = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=A�A�A�A��LD�����3333DDDD    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( �A�LDL�L�D�L�����3333DDDD x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx""""wwwwwwDGAD w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww""""wwwwqqDAAq  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(""""wwwwwwwGGwGGwGwGw �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((�UQUUQUUQUUQUUUDUUUUU3333DDDD ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`DEQQUUDUTEUUUU3333DDDD M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M""""������������������������ � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""�������DAADAI � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(��A�AM�M�DM��M334CDDDD 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5DD����M��DM�����3333DDDD x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x""""wwwwwwDGqGq w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwwGwwDGwwwwwwww + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+ADAH�DJ�H�H�����3333DDDD � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(��H��J�AD�DH�D����3333DDDD � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�""""�������DD����� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
� �@kV` k^ �c� � c� � �C. � C6  C7! �	C8! � 
C: � C; �J�
 �J� �J� �J� �J� �C' � C"- �C#  �C%( � C'0 �kj �kr � �c� � �c� � � c� � �	� � �	� � �� � �� � xC � x  C � y !C � q "C � i #C � a $C � �%"� � � &"� � �'"� � �(*� � z )*OW z**(_ �+**o �,*8g � -*Gg � .*Ew � /*Pg �0" �1*o 2*Fg3)�w*4*8g: 5*Gg:  *Ew: 7*Gg:  *Ew: 9*JwJ )�g �;)�g �<**=*<g
>*2w* *:g3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�������������������������������������������=�K�K�S�[��<�K�R�G�T�T�K� � � � � � � �@�9�1����������������������������������������� ��=�K�X�X�_��B�G�Q�K� � � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������@�9�1� ���������������������������������������2�0�.�	�
�������������������� � � � � � �����������������������������������������%��������������������2�0�.� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            