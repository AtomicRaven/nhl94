GST@�                                                           �e�                                                       �� ��U �c�~   ��	         j�������J���ʰ���������    ����        2:     #    ����                                d8<n    �  ?     �����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    "�j��,  " ��
  �                                                                               ����������������������������������      ��    oo? 0 go5  8  +     '        ��  
    
          	� 74 V 	�                 �Y          8::�����������������������������������������������������������������������������������������������������������������������������?o  0  5o  8    +     '            �  
     
            �	  47  V  �	                  Y            :: �����������������������������������������������������������������������������                                         �   @  &   }   �                                                                                 'w w  �Y  Y    �0   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E E �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    L��bD�X&=4m �L3��{�E��qA�P^^��_X13�T0 k� �,{�0{U2d  9U8D"!  ��3    � )�8L��cD�X(=4n �L7��{�E��sA�P^^��_X13�T0 k� �4{�8{U2d  9U8D"!  ��3    � )�8L��dD�\*=8n �L7��{�E� tA�T_^��_T13�T0 k� �<{�@{U2d  9U8D"!  ��3    � )�8L��eD�\,=<n �L;��{�E�vA�T_^��_P13�T0 k� �@{�D{U2d  9U8D"!  ��3    � )�8L��fD�\.=@o  L;��{�E�wA�T_^�_P13�T0 k� �H{�L{U2d  9U8D"!  ��3    � )�8L��gD�\0MDo L?��w�B�yA�X_^�_L13�T0 k� �L{�P{U2d  9U8D"!  ��3    � )�8L��hL|`2MDo L?��{�B�{A�X_^{�_L13�T0 k� �T{�X{U2d  9U8D"!  ��3   � )�8L��iL|`4MHo �LC��{�B�|A�\_^{�_H13�T0 k� �X{�\{U2d  9U8D"!  ��3    � )�8L��jL|`6MLp \C��{�B�}A�\_^w�_H13�T0 k� �`{�d{U2d  9U8D"!  ��3    � )�8L��jL|`8MLp \C��{�B�$~A�`_^w�_D13�T0 k� �d{�h{U2d  9U8D"!  ��3    � )�8L��kL|d:MPp $\G���B�0A�``^s�_D13�T0 k� �l{�p{U2d  9U8D"!  ��3    � )�8L��lL|d;MTp (\G���B�<A�d`^s�_@13�T0 k� �pz�tzU2d  9U8D"!  ��3    � )�8L��mL|d=MTp 0~\K���B�H�A�d`^o�_@13�T0 k� �tz�xzU2d  9U8D"!  ��3    � )�8L��nL|d?MXq 0~\K���B�T�A�d`^o�_<13�T0 k� �|z��zU2d  9U8D"!  ��3    � )�8L��oL|dAM\q 4~\K����B�`�A�h`^o�_<13�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8L��pL|hBM`p 8~\O����B�l�A�h`^k�_<13�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8L��qL|hDMdp <~\O����B�xA�l`^k�_813�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8L��qL|hFMdp -@~\O����B��A�l`^g�_813�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8L��rL|hGMhp -D~\S����B��A�l`^g�_413�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8L��sL|hIMhp -D~lS����B��A�p`^g�_413�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8L��tL�lJMlp -H~lS����B��~A�p`^c�_013�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8L��tL�lLMlp -LlW����B��~A�p`^c�_013�T0 k� ��{��{U2d  9U8D"!  ��3    � )�8L��uL�lMMlp}PlW����B��~A�t`^_�_013�T0 k� ��|��|U2d  9U8D"!  �3    � )�8T��tL�lOMpp}TlW����O��}A�t`^_�_,13�T0 k� ��|��|U2d  9U8D"!  ��3    � )�8T��sL�lPMpp}Xl[����O��}A�t`^_�_,13�T0 k� �|}��}U2d  9U8D"!  ��3    � )�8T��sL�pRMpp}\l[����O��}A�x`^[�_,13�T0 k� �t}�x}U2d  9U8D"!  ��3    � )�8T��rL�pSMtp}`l[����O��|A�x`^[�_(13�T0 k� �p}�t}U2d  9U8D"!  ��3    � )�8T��qL�pUMtp}dl_����O��|A�x`^[�_(13�T0 k� �p}�t}U2d  9U8D"!  ��3    � )�8T��pL�pVMtp}hl_����O��|A�|`^W�_$13�T0 k� �p}�t}U2d  9U8D"!  ��3    � )�8T� oL�pWMxp}ll_����O��{A�|`^W�_$13�T0 k� �p}�t}U2d  9U8D"!  ��3    � )�8T�oL�pYMxp}p|c����O��{A�|`^W�_$13�T0 k� �p}�t}U2d  9U8D"!  ��3    � )�8T�nL�tZMxp}t|c����O��zA��`^S�_ 13�T0 k� �t}�x}U2d  9U8D"!  ��3    � )�8T�mL�t[M|p}x|c����O��zA��`^S�_ 13�T0 k� �x}�|}U2d  9U8D"!  ��3    � )�8T�lL�t]M|p}||c����O��zA��`^S�_ 13�T0 k� �|}��}U2d  9U8D"!  ��3    � )�8T�lL�t^M|p��|g����O��yA��`^O�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�kL�t_M|p��|g����O��yA��`^O�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�jL�t`M|p���|g����O��yA��`^O�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�iL�xbM�p���|k����O��yA��`^K�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�iL�xcM�p���|k����O��xA��`^K�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T� hL�xdM�p���|k����O� xA��`^K�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�$gL�xeM�p���|k����O�xA��`^G�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�(gL�xfM�p���Lo�� ��O�wA��`^G�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�(fL�xgM�p���Lo�� ��O�wA��`^G�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�,eL�|hM�p���Lo�� ��O�wA��`^G�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�0eL�|iM�p���Lo�� ��O�vA��`^C�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�0dL�|jM�p���Ls�� ��O�vA��_^C�_13�T0 k� ��}��}U2d  9U8D"!  ��3   � )�8T�4cL�|l=�p���Ls�� ��O�vA��_^C�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�8cL�|m=�p���Ls�� ��O� vA��_^C�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�8bL�|n=�p���<s�� ��O�$uA��_^?�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�<bL�|o=�p���<w�� ��B�(uA��_^?�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�@aL�|p=�o��<w�� ��B�,uA��_^?�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�@aL��p=�o��<w�� ��B�0uA��_^?�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�D`L��qm�o��<w�� ��B�4tA��_^;�_13�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8T�D_L��rm�o��,{�� ��B�8tA��_^;�_13�T0 k� ��|��|U2d  9U8D"!  ��3    � )�8T�H_L��sm�o��~,{��!��B�DtA��_^;�_13�T0 k� ��|��|U2d  9U8D"!  ��3    � )�8T�L^L��tm�o��~,��!��B�LtA��_^;�_13�T0 k� ��|��|U2d  9U8D"!  ��3    � )�8T�L^L��um�o��~,��!��B�XsA��^^;�_13�T0 k� ��|��|U2d  9U8D"!  ��3    � )�8T�P]L��v]�o��~,��!��B�XsA��^^7�_13�T0 k� ��{��{U2d  9U8D"!  �3   � )�8T�P]L��w]�o��}����!��B�\sA��^^7�_13�T0 k� ��{��{U2d  9U8D"!  ��3    � )�8T�T\L��x]�n��}����!��O`sA��^^7�_13�T0 k� ��{��{U2d  9U8D"!  ��3   � )�8T�X[L��y]�n��}����!��O`sA��^^3�_ 13�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8T�X[L|�z�n��}����!��OdsA��^^3�_ 13�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8T�X[L|�{�n��|����!��OhsA��]^3�_ 13�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8T�X[L|�|�n��|����!��OhsA��]^3�_ 13�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8T�\ZL|�}�m��|����!��OlsA��]^3�^�13�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8T�\ZL|�}�m��|�� �!��OpsA��]^/�^�13�T0 k� ��y��yU2d  9U8D"!  ��3    � )�8T�\ZL|�~-�m��|���!��OtrA��]^/�^�13�T0 k� ��y��yU2d  9U8D"!  ��3    � )�8T�\ZD܄-�l��{���!��OxrA��]^/�^�13�T0 k� ��y��yU2d  9U8D"!  ��3    � )�8T�\ZD܈-�l��{���!��O|rA��\^/�^�13�T0 k� ��y��yU2d  9U8D"!  ��3    � )�8T�\YD܈~-�l��{��"��O�rA��\^/�^�03�T0 k� ��y��yU2d  9U8D"!  ��3    � )�8T�`YD܈~-�k��{�
�"��O�rA��\^/�^�03�T0 k� ��x��xU2d  9U8D"!  ��3    � )�8T�`XD܈~-�k��{��"��O�rA��\^+�^�03�T0 k� ��x��xU2d  9U8D"!  ��3   � )�8T�`XF�~=�j��z��"��O�rA��\^+�^�03�T0 k� ��x��xU2d  9U8D"!  ��3    � )�8T�dXF�}=�j��z��"��O�rA��\^+�^�03�T0 k� ��x��xU2d  9U8D"!  ��3    � )�8T�dWF�}=�j}�z���"��O�rA��[^+�^�03�T0 k� ��x��xU2d  9U8D"!  ��3    � )�8T�dWF�}=�i}�z���"��O�rA��[^+�^�03�T0 k� ��x��xU2d  9U8D"!  ��3    � )�8T�dWF�}=�i}�z���"��O�rA��[^+�^�03�T0 k� ��w��wU2d  9U8D"!  ��3    � )�8T�hVE��|=�i}�z���"��O�qA��[^'�^�03�T0 k� ��w��wU2d  9U8D"!  ��3    � )�8T�hVE��|=�i}�y���"��O�qA��[^'�^�03�T0 k� ��w��wU2d  9U8D"!  ��3    � )�8T�hUE��|=�h}�y���"��O�qA��[^'�^�03�T0 k� ��w��wU2d  9U8D"!  ��3    � )�8T�lUE��|=�h��y���"��O�qA��[^'�^�03�T0 k� ��r��rU2d  9U8D"!  ��3    � )�8T�lUE��{=�h��yL� �"��O�qA��[^'�^�03�T0 k� ��m��mU2d  9U8D"!  ��3    � )�8T�lTE��{=�g��yL�"�"��O�qA��Z^'�^�03�T0 k� ��j� jU2d  9U8D"!  ��3    � )�8T�lTE��{=�g��xL�$�"��B��qA��Z^'�^�03�T0 k� �h�hU2d  9U8D"!  ��3    � )�8T�pTE��{=�g��xL�&�"��B��qA��Z^#�^�03�T0 k� �f�fU2d  9U8D"!  ��3    � )�8T�pSE��z=�f}�xL�(�"��B��qA��Z^#�^�03�T0 k� �c�cU2d  9U8D"!  ��3    � )�8T�pSE��z=�f}�wL�)�"��B��qA��Z^#�^�03�T0 k� �b�bU2d  9U8D"!  ��3    � )�8T�pSE��z=�f}�wL�+�"��B��qA��Z^#�^�03�T0 k� �`�`U2d  9U8D"!  ��3    � )�8T�tRE��y=�f~ vL�-""��@�qA��Z^#�^�03�T0 k� �_�_U2d  9U8D"!  ��3    � )�8T�tRE��y=�e~vL�/"#��@�pA��Z^#�^�03�T0 k� �^�^U2d  9U8D"!  ��3    � )�8T�tRE��x=�euL�1"#��@�pA��Z^#�^�03�T0 k� �^�^U2d  9U8D"!  ��3    � )�8T�tRE��x> euL�3"#��@�pA��Y^#�^�03�T0 k� �^�^U2d  9U8D"!  ��3   � )�8T�xQE��w> duL�5"#��@�pA��Y^�^�0"s�T0 k� �^�^U2d  9U8D"!  ��3    � )�8T�xQE��v>dt\�7"#��@�pA��Y^�^�0"s�T0 k� �^�^U2d  9U8D"!  ��3    � )�8T�xQE��v>dt\�9"#��@�pA��Y^�^�0"s�T0 k� �]�]U2d  9U8D"!  ��3    � )�8T�xPCL�u>c�s\�;"#��@�oA��Y^�^�0"s�T0 k� �^�^U2d  9U8D"!  ��3    � )�8T�xPCL�t>c�s\�="#��@�oA��Y^�^�0"s�T0 k� �_�_U2d  9U8D"!  ��3    � )�8T�|PCL�s>b�s\�?"#��@�oA��Y^�^�0"s�T0 k� �_�_U2d  9U8D"!  ��3   � )�8T�|PCL�r>b� r	\�A"#��@�oA��Y^�^�0"s�T0 k� �_�_U2d  9U8D"!  ��3    � )�8T�|OCL�r>b� r	\�B�#��@�oA��Y^�^�0"s�T0 k� �^�^U2d  9U8D"!  ��3    � )�8T�|OCL�q>a~$q	\�D�#��@�oA��Y^�^�0"s�T0 k� �^�^U2d  9U8D"!  ��3    � )�8T��OCL�p>a~(q	\�E�#��@�oA��X^�^�0"s�T0 k� �]�]U2d  9U8D"!  ��3    � )�8T��OK��o>a~(q	\�G�#��@�nA��X^�^�0"s�T0 k� �]�]U2d  9U8D"!  ��3    � )�8T��NK��n>`~(q��H�#��@�nA��X^�^�03�T0 k� �]�]U2d  9U8D"!  ��3    � )�8T��NK��m>`~,p��J�#��@�nA��X^�^�03�T0 k� �]�]U2d  9U8D"!  ��3   � )�8T��NK��l>`~0p��K�#��@�nA��X^�^�03�T0 k� �]�]U2d  9U8D"!  ��3    � )�8T��NK��k> _~0p��M�#��@�nA��X^�^�03�T0 k� �\�\U2d  9U8D"!  ��3    � )�8T��MK��j> _~4o��N�#��@�nA��X^�^�03�T0 k� �\�\U2d  9U8D"!  ��3    � )�8T��MK��i>$^~4o��P�#��@�nA��X^�^�03�T0 k� �[�[U2d  9U8D"!  ��3   � )�8T��MK��h>$^~8o��Q�#��@�nA��X^�^�03�T0 k� �[� [U2d  9U8D"!  ��3    � )�8T��MK��g>(^�<n��R",#��@�mA��X^�^�03�T0 k� � [�$[U2d  9U8D"!  ��3   � )�8T��MK��g>(^�<n��T",#��@�mA��X^�^�03�T0 k� � Z�$ZU2d  9U8D"!  ��3    � )�8T��LK��f>(]�@m��U",#��@�mA��X^�^�03�T0 k� �$Z�(ZU2d  9U8D"!  ��3    � )�8T��LK��e>,]�@m��V",#��@�mA��X^�^�03�T0 k� �$Z�(ZU2d  9U8D"!  ��3    � )�8T��LK��e>,]�Dm��V",#��@�mA��W^�^�0"��T0 k� �8Y�<YU2d  9U8D"! �3    � )�8T��LK� e>0\�Dl��V",#��@ mA��W^�^�0"��T0 k� �LY�PYU2d  9U8D"! ��?    � )�8T��KK�e>0\�Hl��W",#��@ mA��W^�^�0"��T0 k� �\Y�`YU2d  9U8D"! ��?    � )�8T��KK�e>0\�Ll��W",$��@mA��W^�^�0"��T0 k� �pY�tYU2d  9U8D"! ��?    � )�8T��KK�f>4[�Lk��X",$��@mA��W^�^�0"��T0 k� ��Y��YU2d  9U8D"! ��?    � )�8T��KK�f>4[�Pk��X",$��@lA��W^�^�0"��T0 k� ��X��XU2d  9U8D"! ��?    � )�8T��KK�f>8[�Pk��Y",$��@lA��W^�^�0"��T0 k� ��X��XU2d  9U8D"! ��?    � )�8T��KK�f>8[�Tj��Y�$��@lA��W^�^�0"��T0 k� ��X��XU2d  9U8D"!	 ��?    � )�8T��JK�f>8Z�Tj��Z�$��@lA��W^�^�0"��T0 k� ��X��XU2d  9U8D"!
 ��?   � )�8T��JK�f><Z�Xj��Z�$��@lA��W^�^�0"��T0 k� ��X��XU2d  9U8D"! ��?    � )�8T��JK� f><Z�Xj��[�$��@lA��W^�^�0"��T0 k� ��X��XU2d  9U8D"! ��?    � )�8T��JK�$f><Z�\i��[�$��@lA��W^�^�03�T0 k� �W�WU2d  9U8D"! ��?    � )�8T��JK�(f>@Y�\i��\�$��@lA��W^�^�03�T0 k� �W� WU2d  9U8D"! ��?    � )�8T��JK�,f>@Y�\i��\�$��@lA��W^�^�03�T0 k� �0W�4WU2d  9U8D"! ��?    � )�8T��IK�,f>@Y�`h��]�$��@lA��W^�^�03�T0 k� �@W�DWU2d  9U8D"! ��?    � )�8T��IK�0f>DY�`h��]�$��@lA��W^�^�03�T0 k� �TW�XWU2d  9U8D"! ��?    � )�8T��IK�4f>DX�dh��]�$��@kA��V^�^�03�T0 k� �hV�lVU2d  9U8D"! ��?    � )�8T��IK�8g>DX�dh��^�$��@kA��V^�^�03�T0 k� �xV�|VU2d  9U8D"! ��?    � )�8T��IK�8g>HX�hg��^�$��@kA��V^�^�03�T0 k� ��V��VU2d  9U8D"! ��?    � )�8T��IK�<g>HX�hg��_�$��@kA��V^�^�03�T0 k� ��V��VU2d  9U8D"! ��?    � )�8T��HK�@g>HX�lg��_�$��@ kA��V^�^�03�T0 k� ��V��VU2d  9U8D"! ��?    � )�8T��HK�Dg>LW�lg��_�$��@ kA��V^�^�03�T0 k� ��V��VU2d  9U8D"! ��?    � )�8T��HK�Dg>LW�lf��`�$��@ kA��V^�^�03�T0 k� ��U��UU2d  9U8D"! ��?    � )�8T��HK�Hg>LW�pf��`�$��@$kA��V^�^�03�T0 k� ��U��UU2d  9U8D"! ��?    � )�8U�HK�Lg>PW�pf��a�$��@$kA��V^�^�03�T0 k� � U�UU2d  9U8D"! ��?    � )�8U�HK�Lg>PV�pf��a�$��@$kA��V^�^�03�T0 k� �U�UU2d  9U8D"! ��?    � )�8U�HK�Pg>PV�te��a�$��@(kA��V^�^�03�T0 k� �$U�(UU2d  9U8D"! ��?    � )�8U�GK�Tg>PV�te��b�$��@(kA��V^�^�03�T0 k� �8U�<UU2d  9U8D"! ��?    � )�8U�GK�Tg>TV�xe��b�$��@(kA��V^�^�03�T0 k� �LT�PTU2d  9U8D"! ��?   � )�8U�GK�Xg>TV�xe��b�$��@,jA��V^�^�03�T0 k� �\T�`TU2d  9U8D"! ��?    � )�8U�GK�Xg>TV�xe��c�$��@,jA��V^�^�03�T0 k� �pT�tTU2d  9U8D"! ��?    � )�8U�GK�\g>TU�|d��c�$��@,jA��V^�^�03�T0 k� ��T��TU2d  9U8D"! ��?    � )�8U�GK�`h>XU�|d��c�$��@,jA��V^�^�03�T0 k� �T��TU2d  9U8D"! ��?    � )�8U��GK�`h>XU�|d��d�$��@0jA��V^�^�03�T0 k� �S��SU2d  9U8D"! ��?    � )�8U��GK�dh>XU��d��d�$��@0jA��V^�^�03�T0 k� �S��SU2d  9U8D"! ��?    � )�8U��GK�dh>XU��c��d�$��@0jA��V^�^�03�T0 k� ��S��SU2d  9U8D"! ��?    � )�8U��FK�hh>\T��c��e�$��@4jA��V^�^�03�T0 k� ��S��SU2d  9U8D"! ��?    � )�8U��FK�lh>\T��c��e�$��@4jA��V^�^�03�T0 k� ��S��SU2d  9U8D"! ��?    � )�8U��FK�lh>\T��c��e�$��@4jA��V^�^�03�T0 k� �S�SU2d  9U8D"! ��?    � )�8U��FK�ph>\T��c��e�$��@4jA��V^�^�03�T0 k� �R� RU2d  9U8D"! ��?    � )�8U��FK�ph>`T��c��f�$��@8jA��U^�^�03�T0 k� �,R�0RU2d  9U8D"! ��?    � )�8U��FK�th>`T��b��f�%��@8jA��U^�^�03�T0 k� �@R�DRU2d  9U8D"! ��?    � )�8DݜFK�th>`T��b��f�%��@8jA��U^�^�03�T0 k� �TR�XRU2d  9U8D"! ��?    � )�8DݜFK�xh>`S��b��g�%��@8jA��U^�^�03�T0 k� �hR�lRU2d  9U8D"! ��?    � )�8DݜFK�xh>dS��b��g�%��@<jA��U^�^�03�T0 k� �xR�|RU2d  9U8D"! ��?    � )�8DݜFK�|h>dS��b��g�%��@<iA��U^�^�03�T0 k� �Q��QU2d  9U8D"! ��?    � )�8DݠFK�|h>dS��b��g�%��@<iA��U^�^�03�T0 k� �Q��QU2d  9U8D"! ��?    � )�8L]�FK݀h>dS��a��h�%��@<iA��U^�^�03�T0 k� �Q��QU2d  9U8D"! ��?    � )�8L]�FK݀h>dS��a��h�%��@@iA��U^�^�03�T0 k� ��Q��QU2d  9U8D"! ��?    � )�8L]�FCM�h>hS^�a��h�%��@@iA��U^�^�03�T0 k� ��Q��QU2d  9U8D"! ��?   � )�8L]�FCM�h>hR^�a��h�%��@@iA��U^�^�03�T0 k� ��P��PU2d  9U8D"! ��?    � )�8L]�FCM�h>hR^�a��h�%��@@iA��U^�^�03�T0 k� ��P� PU2d  9U8D"! ��?    � )�8L]�FCM�h>hR^�a��h�%��@DiA��U^�^�03�T0 k� �P�PU2d  9U8D"! ��?    � )�8L]�GCM�h>hR^�`��h�%��@DiA��U^�^�03�T0 k� �$P�(PU2d  9U8D"! ��?    � )�8L]�GCM�g>hR^�`��h�%��@DiA��U^�^�03�T0 k� �8P�<PU2d  9U8D"! ��?    � )�8L]�GE��g>lR^�`�h�%��@DiA��U^�^�03�T0 k� �HP�LPU2d  9U8D"! ��?    � )�8L]�GE��g>lR^�`�h�%��@DiA��U^�^�03�T0 k� �\O�`OU2d  9U8D"! ��?    � )�8L]�GE��f>lR^�`�h�%��@HiA��U^�^�03�T0 k� �pO�tOU2d  9U8D"! ��?    � )�8L]�GE��f>lQ^�`�h�%��@HiA��U^�^�03�T0 k� �O��OU2d  9U8D"! ��?    � )�8L]�GE��eNlQn�`�h�%��@HiA��U^�^�03�T0 k� �O��OU2d  9U8D"! ��?    � )�8Lm�GE͔eNpQn�_�h�%��@HiA��U^�^�03�T0 k� �O��OU2d  9U8D"! ��?    � )�8Lm�GE͔dNpQn�_\�h�%��@HiA��U^�^�03�T0 k� �O��OU2d  9U8D"! ��?    � )�8Lm�GE͘dNpQn�_\�h�%��@LiA��U^�^�03�T0 k� ��N��NU2d  9U8D"! ��?    � )�8Lm�GE͘cNpQn�_\�h�%��@LiA��U^�^�03�T0 k� ��N��NU2d  9U8D"! ��?    � )�8Lm�GE͘bNpQn�_\�h�%��@LiA��U^�^�03�T0 k� ��N��NU2d  9U8D"! ��?    � )�8Lm�GE͘bNpQn�_\�h�%��@LiA��U^�^�03�T0 k� �N�NU2d  9U8D"! ��?    � )�8Lm�GEݘaNtQn�_��h�%��@LiA��U^�^�03�T0 k� �N�NU2d  9U8D"! ��?    � )�8Lm�GEݘ`NtPn�_��h�%��@LiA��U^�^�03�T0 k� �,M�0MU2d  9U8D"! ��?    � )�8Lm�HEݘ`^tP^�_��h�%��@PiA��U^�^�03�T0 k� �@M�DMU2d  9U8D"! ��?    � )�8Lm�HEݘ_^tP^�^��h�%��@PiA��U^�^�03�T0 k� �TM�XMU2d  9U8D"! ��?    � )�8Lm�HEݘ^^tP^�^��h�%��@PhA��U^�^�03�T0 k� �dM�hMU2d  9U8D"! ��?    � )�8Lm�HEݘ^^tP^�^��h�%��@PhA��U^�^�03�T0 k� �xM�|MU2d  9U8D"! ��?    � )�8Lm�HEݘ]^tP^�^��h�%��@PhA��U^�^�03�T0 k� �M��MU2d  9U8D"! ��?    � )�8Lm�HEݔ]^xP^�^��h�%��@PhA��U^�^�03�T0 k� �L��LU2d  9U8D"! ��?    � )�8Lm�HEݔ\^xP^�^��h�%��@ThA��U^�^�03�T0 k� �L��LU2d  9U8D"! ��?    � )�8Lm�HK�[^xP^�^��h�%��@ThA��U^�^�03�T0 k� ��L��LU2d  9U8D"! ��?    � )�8Lm�HK�[^xP^�^��h�%��@ThA��U^�^�03�T0 k� ��L��LU2d  9U8D"! ��?    � )�8Lm�HK�ZxP��^��g�%��@ThA��U^�^�03�T0 k� ��L��LU2d  9U8D"! ��?    � )�8Lm�HK�YxO��]��g�%��@ThA��U^�^�03�T0 k� ��L� LU2d  9U8D"! ��?    � )�8Lm�HK�YxO��]��g�%��@ThA��U^�^�03�T0 k� �K�KU2d  9U8D"! ��?   � )�8Lm�HEm�XxO��]��g�%��@XhA��U^�^�03�T0 k� �$K�(KU2d  9U8D"! ��?    � )�8Lm�HEm�W|O��]��f�%��@XhA��U^�^�03�T0 k� �4K�8KU2d  9U8D"! ��?    � )�8Lm�HEm�V|O��]��f�%��@XhA��U^�^�03�T0 k� �HK�LKU2d  9U8D"! ��?    � )�8Lm�HEm�V|O^�]��f�%��@XhA��U^�^�03�T0 k� �\K�`KU2d  9U8D"! ��?    � )�8Lm�HEm�V|O^�]��f�%��@XhA��U^�^�03�T0 k� �pJ�tJU2d  9U8D"!
 ��?   � )�8C�PC�߇�7���/�|?��3�E�;Ea�	���DS3�T0 k� ��7��7U2d  9U8D"!  ��'    � ��C� PC�׆�+���/�|?��+�E�:EQ�	���HT3�T0 k� ��8��8U2d  9U8D"!  ��'    � ��C��OC�ӆ�#���.�|?��#�E�:EQ�	À�HU3�T0 k� ��9��9U2d  9U8D"!  ��'    � ��C��OC�˅�� �-�|?���E� :EQ�	À�LV3�T0 k� ��>��>U2d  9U8D"!  ��'    � ��C��OC�Å�� �-�|?���E��:EQ�	À�LW3�T0 k� ��B��BU2d  9U8D"!  ��'    � ��C��NC⿄�� �,�|?���E��:EQ�	À�PX3�T0 k� ��E��EU2d  9U8D"!  ��'    � ��C��MC⯃��� �,�|?����E��:C��	���TZ3�T0 k� ��G��GU2d  9U8D"!  ��'    � ��C��LC⧃��� �,��|?����E��;C��	���X[3�T0 k� ��J��JU2d  9U8D"!  ��'    � ��C��LC⟃��� �,��|?����E��;C��	���\\3�T0 k� �K��KU2d  9U8D"!  ��'    � ��C��KC���� �,��|?����E��;C���	��s`\3�T0 k� �L��LU2d  9U8D"!  ��'    � ��C��KC���� �,�||?����A��;C���	��s`]3�T0 k� �K��KU2d  9U8D"!  ��'    � ��C��JC���� �,�x|?����A��<C�����sd]3�T0 k� �K��KU2d  9U8D"!  ��'    � ��C��JC���� �,�p|?����A��<C�����sh^3�T0 k� �J��JU2d  9U8D"!  ��'    � ��C��IC�{�ߴ�+`l|?����A��<C�����sl^3�T0 k� ��I��IU2d  9U8D"!  ��'    � ��C��HC�s�߬x+`h|?����A��=C�����sl_3�T0 k� ��J��JU2d  9U8D"!  ��'    � ��EрHC�k�ߨt+``|?���A��=C�����sp_3�T0 k� �|J��JU2d  9U8D"!  ��'    � ��E�xGC�c�ߠl+`\|?���A��>C�����st_3�T0 k� �tK�xKU2d  9U8D"!  ��'    � ��E�hFC�S�ߐ\+`P|?���A��?C������x`3�T0 k� �hL�lLU2d  9U8D"!  ��'    � ��E�`FC�K�߈	T+`L|?���A��?EP��S��|`3�T0 k� �`L�dLU2d  9U8D"!  ��'    � ��E�XEDC�߀
L+`D|?���A��@EP��S��|`3�T0 k� �XM�\MU2d  9U8D"!  ��'    � ��E�PED;��xD*`@|?���A��AEP��S���`3�T0 k� �PN�TNU2d  9U8D"!  ��'    � ��C�HDD3��p<*`8|?���A�xAEP��S���`3�T0 k� �HN�LNU2d  9U8D"!  ��'    � ��C�@DD+��l4*`4|?���A�pBEP��S���`3�T0 k� �@O�DOU2d  9U8D"!  ��'    � ��C�4CD#��d�,*`,|?��w�A�hCEP��S���`3�T0 k� �8P�<PU2d  9U8D"!  ��'    � ��C�,CD��\�$*P$|?�1o�A�`DEP� S���`3�T0 k� �0Q�4QU2d  9U8D"!  ��'    � ��C�$BD��T�*P |?�1g�A�XEEP� S���_3�T0 k� �(R�,RU2d  9U8D"!  ��'    � ��E�BD��L�*P|?�1c�EPPEE@�S���_3�T0 k� �$L�(LU2d  9U8D"!  ��'    � ��E�AD��D�*P|?�1[�EPHFE@�S���_3�T0 k� � I�$IU2d  9U8D"!  ��'    � ��E�AD���@�*P|?�1S�EP@GE@�S���_3�T0 k� �G�GU2d  9U8D"!  ��'    � ��E�@D��8��*P|?�1K�EP8GE@�S���_3�T0 k� �D�DU2d  9U8D"!  ��'    � ��E��@D�_0��)_�
|?�1C�EP0HE@�S���_3�T0 k� �C�CU2d  9U8D"!  ��'    �  ��E��@D�_(��)_�	|?�1;�EP(IE@�S���_3�T0 k� �C�CU2d  9U8D"!  ��'    � !��E��?Dۅ_$��)��|?�17�EP IE@|S���_3�T0 k� ��C� CU2d  9U8D"!  ��'    � !��E��?DӅ_��)��|?�1/�EPJE@xS���_3�T0 k� ��B��BU2d  9U8D"!  ��'    � "��E��>Dυ_��)��|?�1'�EPKE@pS���_3�T0 k� ��B��BU2d  9U8D"!  ��'    � #��E��>Dǅ_��)��|?�1�EPKC�hS���_3�T0 k� ��B��BU2d  9U8D"!  ��'    � #��E��>D��_��(��|?�A�E_�LC�dS���_3�T0 k� ��C��CU2d  9U8D"!  ��'    � $��E�=D��_�(��|?�A�E_�MC�\S���_3�T0 k� ��D��DU2d  9U8D"!  ��'    � %��EP�=D��^��(��|?�A�EO�MC�TS���_3�T0 k� ��A��AU2d  9U8D"!  ��'    � %��EP�=D��^��'�|< A�EO�NC�PS���^3�T0 k� ��@��@U2d  9U8D"!  ��'    � &��EP�<D��^�!�'�|8 @��EO�OC�@S���^3�T0 k� ��@��@U2d  9U8D"!  ��'    � '��EP�<CᏆ^�"�&�|8@��EO�OC�<S���^3�T0 k� ��?��?U2d  9U8D"!  ��'    � '��EP�<Cᇇ^�#�&�|8@��EO�OC�4S���^3�T0 k� ��?��?U2d  9U8D"!  ��'    � '��EP�;C��^�$��&�� |8@��A�PC�,S���^3�T0 k� ��?��?U2d  9U8D"!  ��'    � (��C�x;C�w�^�%�|%�� |8@��A�PC�$S���^3�T0 k� ��?��?U2d  9U8D"!  ��'    � (��C�p;C�o�^�%�t%���|8@��A�PC�S���^3�T0 k� �p?�t?U2d  9U8D"!  ��'    � (��C�h:C�g�^�&�l$��|8P��A�QC� S���^3�T0 k� �d?�h?U2d  9U8D"!  ��'    � )��C�`:C�_�^�'�h#�w�|8P��A�QC� S���^3�T0 k� �X?�\?U2d  9U8D"!  ��'    � )��C�T:C�W�^�(�`#�o�|8P��A�QC� S���^3�T0 k� �L?�P?U2d  9U8D"!  ��'    � )��C�L:C�O�^�)�X"�g�|8P��A�QC��S���^3�T0 k� �D?�H?U2d  9U8D"!  ��'    � )��C�D9C�G�^�)�P!�_�|8P��AxQC���S���^3�T0 k� �<?�@?U2d  9U8D"!  ��'    � )��C�<9C�?�^�*�L �W�|8P��AlQC���S���^3�T0 k� �0?�4?U2d  9U8D"!  ��'    � )��C�49C�7�^�+�D �O�|8P��AdQC���S���^3�T0 k� �(?�,?U2d  9U8D"!  ��'    � )��C�,9C�/�^�,�<�G�|8P��A\QC���S���^3�T0 k� � ?�$?U2d  9U8D"!  ��'    � )��C� 8C�'�^�,�8?�|8P��APQC���S���^3�T0 k� �?�?U2d  9U8D"!  ��'    � )��C�8C��^�-�07�|8P��A/HQC���S���^3�T0 k� �?�?U2d  9U8D"!  ��'    � )��C�8C��^�.o(/�|8P��A/@PC���S���^3�T0 k� �?�?U2d  9U8D"!  ��'    � )�C�8C��^�.o$'�|8`�A/4PC���S���^3�T0 k� �>�>U2d  9U8D"!  ��'    � )�}C� 7C��^�/o�|8`w�A/,PC���S���]3�T0 k� ��>��>U2d  9U8D"!  ��'    � )�zC��7C���^�0o�|8`s�A/$PC���S���]3�T0 k� ��>��>U2d  9U8D"!  ��'    � )�xC��7C���^�1o�|8`k�E�PC���S���]3�T0 k� ��C��CU2d  9U8D"!  ��'    � )�vC��7C��^�1o�|8`c�E�PC���S���]3�T0 k� ��F��FU2d  9U8D"!  ��'    � )�sC��6C��^|2n���|8`W�E� OEO��S���]3�T0 k� ��H��HU2d  9U8D"!  ��'    � )�pC��6D ۊ^x3n���|8`O�E��OEO��S���]3�T0 k� ��I��IU2d  9U8D"!  ��'    � )�mC��6D ӊ^t4n���|8`K�E��OEO��S���]3�T0 k� ��K��KU2d  9U8D"!  ��'    � )�kC��6D ˊ^p4n���|8`C�E��OEO��S���]3�T0 k� ��L��LU2d  9U8D"!  ��'    � )�hD�5D Ê^l5^���|8`;�An�OEO�S���]3�T0 k� ��L��LU2d  9U8D"!  ��'    � )�fD�5D ��^h6^���|807�An�OEOw�S���]3�T0 k� ��L��LU2d  9U8D"!  ��'    � )�dD�5D ��^d6^���|80/�An�NEOo�S���]3�T0 k� ��L��LU2d  9U8D"!  ��'    � )�aD�5D ��^`7^���|80'�An�NEOg�S���]3�T0 k� �tK�xKU2d  9U8D"!  ��'    � )�_D�5D ��^\7^���|80#�An�NEO_�S���]3�T0 k� �hK�lKU2d  9U8D"!  ��'    � )�\D�5D ��^X8^���|80�E^�NEO[����]3�T0 k� �lI�pIU2d  9U8D"!  ��'    � )�ZD|4D ���T8^�
��|80�E^�NE?S����]3�T0 k� �lH�pHU2d  9U8D"!  ��'    � )�XDl4D ���L9^���|80�E^�NE?C����\3�T0 k� �`G�dGU2d  9U8D"!  ��'    � )�VD`4D{��H:^���|80�E^�NE??����\3�T0 k� �\F�`FU2d  9U8D"!  ��'    � )�TDX4Ds��D:^���|8?��EN�ME?7��|s�\3�T0 k� �TC�XCU2d  9U8D"!  ��'    � )�RDP3Dk��@:N���|8?�ENxME?/��|s�[3�T0 k� �P@�T@U2d  9U8D"!  ��'    � )�PDH3Dc��<;N��{�|8?�ENlME?+��|s�[3�T0 k� �H>�L>U2d  9U8D"!  ��'    � )�ND83DS��4;N|�k�|4O�EN\LE?��xs�Z3�T0 k� �8<�<<U2d  9U8D"!  ��' 
   � )�LD,3DK��0;Nt�c�|4OۺATLE?��tc�Z3�T0 k� �(;�,;U2d  9U8D"!  ��' 
   � )�JD$3DC��(;Nl�[�|4OӹAHLE?��tc�Y3�T0 k� �;� ;U2d  9U8D"!  ��' 
   � )�HD2D;��$;Nd�S�|4	OϸA@KE?��pc�X3�T0 k� �:�:U2d  9U8D"!  ��' 
   � )�GD2D3�� <N\ �K�|4	OǷA8KE/��lc�X3�T0 k� � :�:U2d  9U8D"!  ��' 
   � )�FD2D+��<�T �C�|4	_��A8KE.���lc�W3�T0 k� ��:��:U2d  9U8D"!  ��' 
   � )�ED�2C���;�K��3�|4	_��A8KE.���dS�V3�T0 k� ��:��:U2d  9U8D"!  ��' 
   � )�DC��2C���;�C��+�|4	_��A0KE.���`S�V3�T0 k� ��9��9U2d  9U8D"!  ��' 
   � )�CC��2C���:�;����4	_��A(KI>���\S�U3�T0 k� ��9��9U2d  9U8D"!  ��' 
   � )�BC��1C���:�3����4	_��A. KI>���XS�U3�T0 k� ��9��9U2d  9U8D"!  ��' 
   � )�AC��1C�����:�+����0	_��A.KI>���TS�T3�T0 k� ��9��9U2d  9U8D"!  ��' 
   � )�@C��1C����9�#����0	_��A.KI>���PS�T3�T0 k� ��9��9U2d  9U8D"!  ��' 
   � )�?C��1C����9������0	_��A.JI>���LS�S3�T0 k� ��8��8U2d  9U8D"!  ��' 
   � )�>C�1C�ߍ��8��]���0
��A-�JIN��D��R3�T0 k� ��8��8U2d  9U8D"!  ��' 
   � )�=C�1C�׍��8��]���0
�w�A-�IIN��@��R3�T0 k� ��7��7U2d  9U8D"!  ��' 
   � )�<C�1C�ύ��8���]���0
�s�A-�IIN��<��Q3�T0 k� ��7��7U2d  9U8D"!  ��' 
   � )�;C�0C�Ǎ��7���]���0
�k�A-�HIN��4��Q3�T0 k� ��7��7U2d  9U8D"!  ��' 
   � )�:C�0C�����7���]���0
�c�A-�HIN��0��P3�T0 k� ��6��6U2d  9U8D"!  ��' 
   � )�9C��0C���m�7���]���0
�[�A-�GI>��,��P3�T0 k� ��5��5U2d  9U8D"!  ��' 
   � )�8C�x0C���m�6���]���0
�O�A=�FI>�� ��O3�T0 k� ��3��3U2d  9U8D"!  ��' 
   � )�8C�l0C���m�6���]���0
�G�A=�FI>���N3�T0 k� �|3��3U2d  9U8D"!  ��' 
   � )�8C�d0C���m�5���]���0�?�A=�EI>���N3�T0 k� �t2�x2U2d  9U8D"!  ��' 
   � )�8C�\0C���m�5���]���0�;�A=�EIN���N3�T0 k� �l2�p2U2d  9U8D"!  ��' 	   � )�8C�T/C���m�4���M���0�3�A=�DIN���M3�T0 k� �d1�h1U2d  9U8D"!  ��' 	   � )�8C�D/C�w�m�3���M���0�#�EM�CIN����L3�T0 k� �T0�X0U2d  9U8D"!  ��' 	   � )�8C�8/C�o�m�2���M��0��EMxBIN����L3�T0 k� �P/�T/U2d  9U8D"!  ��' 	   � )�8C�0/Dg�]�2���Mw��0��EMpAI>����L3�T0 k� �L.�P.U2d  9U8D"!  ��' 	   � )�8D(/D_�]�1���Mo��0��EMhAI>����K3�T0 k� �D.�H.U2d  9U8D"!  ��' 	   � )�8D /DW�]�0�� Mg��0��EM`@I>����K3�T0 k� �<-�@-U2d  9U8D"!  ��' 	   � )�8D/DG�]�/�p MS��0���EMP>I>����J3�T0 k� �,+�0+U2d  9U8D"!  ��' 	   � )�8D.D?�]�.�hMK��0��E=D>@�����J3�T0 k� �,*�0*U2d  9U8D"!  ��' 	   � )�8D�.D7�]�.�`MC��0��E=<=@������|I3�T0 k� �()�,)U2d  9U8D"!  ��' 	   � )�8I��.D/�]|-�XM;��0��E=4<@������tI3�T0 k� � (�$(U2d  9U8D"!  ��' 	   � )�8I��.D'�]t-�P=3��0ۜE=,;@����pI3�T0 k� �'� 'U2d  9U8D"!  ��'    � )�8I��.D�]p,�H=+��0כE=$:@����hH3�T0 k� �&�&U2d  9U8D"!  ��'    � )�8I��.D�]d+�8=��0ǚE=8EΟ��\H3�T0 k� �#�#U2d  9U8D"!  ��'    � )�8I��.D�]\*�0=��0��E=6EΟ��TG3�T0 k� � "�"U2d  9U8D"!  ��'    � )�8I��.D�]T*�(=��0��E�5EΛ��PG3�T0 k� ��"��"U2d  9U8D"!  ��'    � )�8I��.D��]P)� =��0��E��4EΛ��HG3�T0 k� ��"��"U2d  9U8D"!  ��'    � )�8I��.D�]H)�L���0��E��3EΗ��@F3�T0 k� ��"��"U2d  9U8D"!  ��'    � )�8I��.D�]@(�L���0��E��2Eޓ��x8F3�T0 k� ��!��!U2d  9U8D"!  ��'    � )�8I��.Dۏ]4'� L���0��E��/Eޏ��h,E3�T0 k� ����U2d  9U8D"!  ��'    � )�8E]�.DӏM,'��L���0��E��.Eދ��\$E3�T0 k� ����U2d  9U8D"!  ��'    � )�8E]�.DˏM$&�����0��E��-Eދ��TE3�T0 k� ����U2d  9U8D"!  ��'    � )�8E]�.DˏM&l����0�E��,E���LD3�T0 k� ����U2d  9U8D"!  ��'    � )�8E]�.D��M&l����0o�E̸)E���<D3�T0 k� ����U2d  9U8D"!  ��7    � )�8E]�.CM%l����0g�Ḛ(E�{��4�D3�T0 k� ����U2d  9U8D"!  ��7    � )�8E]x.CM %l�ܯ��0
_�Ę&E�w��,�C3�T0 k� ����U2d  9U8D"!  ��7    � )�8E]p.CL�%\�ܧ��0
W�E̠%E�s��$�C3�T0 k� ����U2d  9U8D"!  ��7    � )�8E]l.CL�%\�ܟ��0	O�E̜$E�s���C3�T0 k� ����U2d  9U8D"!  ��7    � )�8E]\.CL�%\�ܓ��0C�E܌!E�k���B3�T0 k� �p�tU2d  9U8D"!  ��7    � )�8E]T.CL�%\�	����0�;�E܄ D>g� ��B3�T0 k� �h�lU2d  9U8D"!  ��7    � )�8EML.CL�%\�	����0�3�E�|D>_����B3�T0 k� �`�dU2d  9U8D"!  ��7    � )�8EMD.CL�%\�	���0�+�E�tD>[���A3�T0 k� �X�\U2d  9U8D"!  ��7    � )�8EM<.C��L�&\�	�w��0�#�E�lD>W���A3�T0 k� �P�TU2d  9U8D"!  ��7    � )�8EM,.C�o�L�&�x	�k��0��G�\D>O���A3�T0 k� �<�@U2d  9U8D"!  ��7    � )�8EM$.E�g�<�&�p	�g��0��G�TD>K���@3�T0 k� �0�4U2d  9U8D"!  �7    � )�8EM-E�_�<�'�p	�_��,��G�PD>G���@3�T0 k� �$�(U2d  9U8D"!  ��3    � )�8EM-E�W�<�'�l	�_��(���G�HD>C���@3�T0 k� � �$U2d  9U8D"!  ��3    � )�8EM,E�K�<�(�d\_��(��G�8E�7���|?3�T0 k� ��U2d  9U8D"!  $�3    � )�8EL�,I�C�<�)�`\[�$��G�0E�3���t?3�T0 k� ,�U2d  9U8D"!  ��?    � )�8EL�,I�;�<x)�`\W�$�ߌG�0E�/���l?3�T0 k� ,�U2d  9U8D"!  ��?    � )�8E<�+I�3�t*�\\S� �׌G�0E�'���d?3�T0 k� ,�U2d  9U8D"!  ��?    � )�8E<�*I�'�d+�\	�O��ˋG�0E����T>3�T0 k� ,�U2d  9U8D"!  ��?    � )�8E<�)I�#�\,�X
�K��ËG�0E��|�L>3�T0 k� ��U2d  9U8D"!  ��?    � )�8E<�)I��T-�X
�G����G�,En�p�D>3�T0 k� ��U2d  9U8D"!  ��?    � )�8E<�(I���L.�T�C����G�,En�h�<>3�T0 k� ��U2d  9U8D"!  ��?    � )�8E<�'I���D/�T�?����G�,En�`�4=3�T0 k� ��U2d  9U8D"!  ��?    � )�8E<�&I���40�T�3����G�,Em��P�$=3�T0 k� ��U2d  9U8D"!  ��?    � )�8E<�%I���,1�T�/�, ���G�,Em���H�=3�T0 k� ��U2d  9U8D"!  ��?    � )�8E<�$I���	�$2�P�+�, ��G�(Em���@=3�T0 k� ��U2d  9U8D"!  ��7    � )�8E<�#I���	�3�P�'�, ��G�(E]���8<3�T0 k� ��� U2d  9U8D"!  ��7    � )�8E<�!I��	�4LL��,  w�G�(E]���$�<3�T0 k� ����U2d  9U8D"!  ��7    � )�8E,� I��	�5LL��,  o�G�(E]����<"��T0 k� ����U2d  9U8D"!  ��7    � )�8E,|I��	� 5LH��+� ]g�G�$E]����<"��T0 k� ����U2d  9U8D"!  ��7    � )�8E,xI��	��6LH��+� ]c�G�$ I�����<"��T0 k� ����U2d  9U8D"!  ��7    � )�8E,xI�ߎ	��7L@��,  ]S�E�$!I������;"��T0 k� ����U2d  9U8D"!  ��7    � )�8E,tI�ێ	��7L8���,  ]K�E�$"I������;"��T0 k� ����U2d  9U8D"!  ��7    � )�8E,pI�ێ	��7L4���,  ]C�E�$"I������;"��T0 k� ����U2d  9U8D"!  ��7    � )�8E,lI�ӎ	��8L,���, ]3�E� $E�����;"��T0 k� ��!��!U2d  9U8D"!  ��7 	   � )�8E,lI�ώ	��8�(���, ]+�G� $E�����:"��T0 k� ��!��!U2d  9U8D"!  ��7 	   � )�8EhE�ώ	��9� ���, ]'�G� %E�����:"��T0 k� �� �� U2d  9U8D"!  ��7 	   � )�8EhE�ˎ	��9����, ]�G�%E�����:3�T0 k� ����U2d  9U8D"!  �7 	   � )�8EdE�Î	��9����, ]�G�&E����:3�T0 k� ����U2d  9U8D"!  ��3 	   � )�8EdEݿ�	��9���, M�G�'E����:3�T0 k� ����U2d  9U8D"!  ��3 	   � )�8B�dE�	��9��, L��G�(E�{���93�T0 k� ����U2d  9U8D"!  ��3 	   � )�8B�`E�	��: ��, L��G�(E�w�0�x93�T0 k� �� �� U2d  9U8D"!  ��3 	   � )�8B�`E�	��:���, L�G�)E�o�0�p93�T0 k� ��"��"U2d  9U8D"!  ��3 	   � )�8B�`E�K�:K���, L߃G�*E�c�0|�`93�T0 k� ��$��$U2d  9U8D"!  ��3 	   � )�8B�`Em��K�:K���, LۃG�*E�[�0t�X93�T0 k� ��%��%U2d  9U8D"!  ��3 	   � )�8B�dEm��K�;K���, LӃG�+E�W�Pl�P93�T0 k� ��&��&U2d  9U8D"!  ��3 	   � )�8B�dEm��K�;K���, L˃G�+E�O�Pd�H8"s�T0 k� ��&��&U2d  9U8D"!  ��3 	   � )�8B�dEm��K�;K���, LÃG�,E�K�P\�@8"s�T0 k� ��'��'U2d  9U8D"!  ��3 
   � )�8B�dE틐K�<K���, L��G�,E�?�PL �08"s�T0 k� ��)��)U2d  9U8D"!  ��3 
   � )�8B�hE퇑K�<K���, L��G�-E�7�PD �(8"s�T0 k� ��*��*U2d  9U8D"!  ��3 
   � )�8B�hE탑K|=K���, L��G�-E�3�P< � 8"s�T0 k� ��+��+U2d  9U8D"!  ��3 
   � )�8B�lE�{�Kt>K����� L��G�.E�+�P7��8"s�T0 k� ��,��,U2d  9U8D"!  ��3 
   � )�8B�lE�w�Kx>K����� L��G�.E�'�P/��8"s�T0 k� ��-��-U2d  9U8D"!  ��3 
   � )�8B�pE�s�Kx>K����� L��G�/F#�P'��7"s�T0 k� ��.��.U2d  9U8D"!  ��3 
   � )�8B�tE�g�K|?K�!������G�0F ����7"s�T0 k� ��0��0U2d  9U8D"!  ��3    � )�8B�xE�c�K|?K�"�����w�G�0F����73�T0 k� ��2��2U2d  9U8D"!  ��3    � )�8B�xE�[�K|@;�#�����o�G�0F����73�T0 k� ��4��4U2d  9U8D"!  ��3    � )�8B�|E�W�K�@;�%�����k�G�1P������73�T0 k� ��6��6U2d  9U8D"!  �3    � )�8E�E�O�;�A;�&�����c�A\1P� �����73�T0 k� ��7��7U2d  9U8D"!  �3    � )�8E�E�G�;�B;�)����S�A\2P��	���P�63�T0 k� ��:��:U2d  9U8D"!  $�3    � )�8E�E�?�;�C;�*����K�A\2P��
	���P�63�T0 k� +�;��;U2d  9U8D"!  ��3    � )�8E�E�;�;�D;�+����G�A\3Q�	���P�63�T0 k� +|=��=U2d  9U8D"!  ��3    � )�8E�E�7�;�D;|-����?�A\3Q�	���P�63�T0 k� +t>�x>U2d  9U8D"!  ��3    � )�8E�E�3�;�E;x.����7�A\4Q�	���P�63�T0 k� +p@�t@U2d  9U8D"!  ��3    � )�8E��D�+�+�F;t0����/�A\4Q�	���P�63�T0 k� +lA�pAU2d  9U8D"!  *�3    � )�8E��D�'�+�G;p1����+�A\ 4Q�	���P�63�T0 k� �lC�pCU2d  9U8D"!  *�3    � )�8E��D�#�+�H;l3����#�A\ 5Q�	���P�63�T0 k� �lD�pDU2d  9U8D"!  *�3    � )�8E��D��+�I �d5�����A\ 5Q�	���P�63�T0 k� �hG�lGU2d  9U8D"!  ��3    � )�8E��D��+�J �h6�����A\ 5Q�	���P�63�T0 k� �dI�hIU2d  9U8D"!  ��3    � )�8BL�D��+�L �h:�����A\ 6P��_��P|53�T0 k� +dL�hLU2d  9U8D"!  ��3    � )�8BL�D��+�M �l;����	�A[�6P��_��Pt53�T0 k� +`N�dNU2d  9U8D"!  ��3    � )�8BL�D��+�N+l=�î�	��A[�7P��_��Pp53�T0 k� +hN�lNU2d  9U8D"!  ��3    � )�8BL�D���O+l?�ì�
��A[�7P��_��Ph53�T0 k� +pO�tOU2d  9U8D"!  ��3    � )�8BL�D����P+pA�ë�
�A[�7P��_��P`53�T0 k� +tO�xOU2d  9U8D"!  ��3    � )�8D��D����Q+pC�Ǫ�
�A[�8D��_�P\53�T0 k� �xQ�|QU2d  9U8D"!  $�3    � )�8D��D����R+pE�ǩ��A[�8D��_{�PT53�T0 k� �xQ�|QU2d  9U8D"!  ��3    � )�8D��D���S+tF�˨��A[�8D��_s�PP53�T0 k� �|S��SU2d  9U8D"!  ��3    � )�8D��D���T {tH�˧�ۋA[�9D��_o�PL53�T0 k� ��W��WU2d  9U8D"!  ��3    � )�8D��D���U {tH�Ϧ�یA[�9D��_k�PD53�T0 k� ��Z��ZU2d  9U8D"!  ��3    � )�8D��D����W {tJ�ϥ�׍A[�9D��_c�P@53�T0 k� ��]��]U2d  9U8D"!  ��3    � )�8D��D����X {xL�Ӥ�ӎA[�9D��__�P843�T0 k� ��_��_U2d  9U8D"!  ��3    � )�8D��D�۷��Z {|O�Ӣ�ˏA[�:D�� _S�P043�T0 k� ��c��cU2d  9U8D"!  ��3    � )�8D��D�׹��[ {�Q�ס�ǐA[�:D��!_O�P(43�T0 k� ��e��eU2d  9U8D"!  ��3    � )�8D��D�ӻ��\+�S�ס�ǑA[�;E|�"_K�P$43�T0 k� ��e��eU2d  9U8D"!  ��3    � )�8D��D�Ͻ��]+�T�ס�ÑA[�;E|�#_G�P 43�T0 k� ��e��eU2d  9U8D"!  ��3    � )�8D��D�Ͼ��^+�V�נ���A[�;E|�$_?�P43�T0 k� ��f��fU2d  9U8D"!  ��3    � )�8D��D�����_+�X�۠���A[�;E|�&_;�P43�T0 k� ��g��gU2d  9U8D"!  ��3    � )�8D��D�����`+�Z�۠���A[�<E} '_7�P43�T0 k� ��h��hU2d  9U8D"!  ��3    � )�8D��D�����b+�^�ߟ���A[�<E}*_/�P43�T0 k� ��l��lU2d  9U8D"!  ��3    � )�8D��D�����c+�`�����A[�<E}+_'�P 43�T0 k� ��m��mU2d  9U8D"!  ��3    � )�8D��D�����d+�a�����A[�=E},_#�_�43�T0 k� ��o��oU2d  9U8D"!  ��3    � )�8D�� D�����e+�c�����A[�=E}._�_�43�T0 k� ��p��pU2d  9U8D"!  ��3    � )�8D��!D�����f+�e�����A[�=D�/_�_�33�T0 k� ��q��qU2d  9U8D"!  ��3    � )�8D��#D���� g�g�����A[�=D�1_�_�33�T0 k� ��m��mU2d  9U8D"!  ��3    � )�8D��%D���h�j�����A��>D�4_�_�33�T0 k� ��m��mU2d  9U8D"!  ��3    � )�8D��&D���i�l�����A��>D�5_�_�33�T0 k� ��l��lU2d  9U8D"!  ��3   � )�8D��(D��� j�m�����A��?A�7_�_�33�T0 k� ��k��kU2d  9U8D"!  ��3    � )�8D��)D���$k�o�����A��?A�8_�_�33�T0 k� ��k��kU2d  9U8D"!  ��3    � )�8D��*D���,l�p�����A��@A�9^��_�33�T0 k� ��k��kU2d  9U8D"!  ��3    � )�8D��,D���4m�q������E��@A�;^��_�33�T0 k� ��l��lU2d  9U8D"!  ��3    � )�8D��-D����<m�r������E��AA�<^��_�33�T0 k� ��l��lU2d  9U8D"!  ��3    � )�8F�/D����Dn +�s������E��AA�=^��_�33�T0 k� ��n��nU2d  9U8D"!  ��3    � )�8F�2D����To +�v������E��CA�@^��_�33�T0 k� �q�qU2d  9U8D"!  ��3    � )�8F�3D����\p +�w������E��CA� A^��_�33�T0 k� �$s�(sU2d  9U8D"!  ��3    � )�8F�5D����dp +�x������E��DA� B^��_�33�T0 k� �0t�4tU2d  9U8D"!  ��3   � )�8F�6D����lq�y�����E��EA�$C^��_�33�T0 k� �,t�0tU2d  9U8D"!  ��3    � )�8F�8D����tq�z�����F�FA�$E^��_�33�T0 k� �(t�,tU2d  9U8D"!  ��3    � )�8F�9D����|r{�����F�GA�$F^��_�33�T0 k� �$u�(uU2d  9U8D"!  ��3    � )�8F�;D�����r|�����F�HA�(G^��_�33�T0 k� �(v�,vU2d  9U8D"!  ��3    � )�8F�=D����r|�����F�IA�(H^��_�23�T0 k� �,v�0vU2d  9U8D"!  ��3    � )�8L|�>D�{���s}�����F�JA�(I^��_�23�T0 k� �0w�4wU2d  9U8D"!  ��3    � )�8L|�@D�{�|�s }�����E{�KA�,J^��_�23�T0 k� �4w�8wU2d  9U8D"!  ��3    � )�8L|�AE�w�|�s�(~�����E{�LA�,K^��_�23�T0 k� �<s�@sU2d  9U8D"!  ��3    � )�8L|�CE�w�|�s�0~�����E{�MA�,M^��_�23�T0 k� �Dq�HqU2d  9U8D"!  ��3    � )�8L|�FE�s�|�s�@~�����E{�PA�0O^��_�23�T0 k� �Xn�\nU2d  9U8D"!  ��3    � )�8L|�GE�o�|�s�H~�����F�QA�0P^��_�23�T0 k� �`l�dlU2d  9U8D"!  ��3    � )�8L|�IE�k�|�s\P�����F�SA�4Q^��_�23�T0 k� �hm�lmU2d  9U8D"!  ��3    � )�8L|�JE�h|�r\X�����F�TA�4R^��_�23�T0 k� �pm�tmU2d  9U8D"!  ��3    � )�8L|�LE�d|�r\`�����F�UA�4S^��_�23�T0 k� �xn�|nU2d  9U8D"!  ��3    � )�8L|�ME�d|�r\h�����F�WA�8T^��_�23�T0 k� ��n��nU2d  9U8D"!  ��3    � )�8L|�NF`|�q\p�����F�XA�8U^��_�23�T0 k� ��n��nU2d  9U8D"!  ��3    � )�8L|�PF`	l�q�x�����F�YA�8V^��_�23�T0 k� ��r��rU2d  9U8D"!  ��3    � )�8L|�QF`l�p�������F�[A�8V^��_|23�T0 k� ��u��uU2d  9U8D"!  ��3    � )�8L��RF\m p�������F�\A�<W^��_x23�T0 k� ��w��wU2d  9U8D"!  ��3    � )�8L��TF\mo�������F�^A�<X^��_x23�T0 k� ��y��yU2d  9U8D"!  ��3    � )�8L��UD�\mo�������D��_A�<Y^��_t23�T0 k� ��z��zU2d  9U8D"!  ��3    � )�8L��VD�\mn�������D��aA�@Z^��_p23�T0 k� ��{��{U2d  9U8D"!  ��3    � )�8L��WD�X=m���#����D��bA�@[^��_p23�T0 k� ��|��|U2d  9U8D"!  ��3    � )�8L��YD�X=m���'����D��dA�@\^��_l23�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8L��ZD�X= l���'����D��fA�@]^��_h23�T0 k� ��}��}U2d  9U8D"!  ��3    � )�8L��[D�X=$l ��+���F�gA�D]^��_h23�T0 k� ��|��|U2d  9U8D"!  ��3    � )�8L��\D�X=$l ��+���F�iA�D^^��_d23�T0 k� ��{��{U2d  9U8D"!  ��3    � )�8L��]D�X=$l ��/���F�jA�H^^��_`23�T0 k� � {�{U2d  9U8D"!  ��3    � )�8L��^D�X =(m ��/���F�lA�H^^��_`23�T0 k� �{�{U2d  9U8D"!  ��3    � )�8L��_D�X"=,m �L3���F�nA�L^^��_\23�T0 k� �{�{U2d  9U8D"!  ��3    � )�8L��aD�X$=0m �L3��{�F�oA�L^^��_\13�T0 k� �${�({U2d  9U8D"!  ��3    � )�8                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��K� ]�#�#� � � H��  � �	    ��l�     H���l��    ��,              
 Z�8           H��    ���   8
           U��  W V
    ��cd?     V>�c�h    ���g              P Z�8          :b  �  ��� 0
% 
           O��   � �       ��k_     O���M(    ���            I Z�8          � �     ���   0
           ]j�   � �
     ����     ]�����    ��Z              j  Z�8          � �     ���  8          f�{   I I   .�7y�     fʗ�7y�                       @	 Z�8          0�  	  ���  P	          %��  ��      B���     %� ���     &                        �             �  ���   P             ��m�          V���    ��g#�     c P              �        �     ��@   09          h��       j����     h�-��r�    ��                  �8          ��     ��J   8�           U �         ~�v�D     Us�v��    �� �                � �         �     ��@   	@
          ����          ���3    ������7      ��               		  ��         	 ��     ��@   H	$
          0��         ���h�     0����m.      ��                A��         
 �     ��@   H
	!          �O ��     � ��9     �O ��9                              ���J             �  ��@      0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          J�  ��        �&� 
@� K�j� >P�UGI�                 x                j  �  �   �                          J    ��        �       K             "                                                �                         �l�c�����7������v���� ���   	 
             
  B   (a� �H�I       / `e� /� f� /� f� 0 f� �d  d@ �  d� ̄ 0\` �� \� � 0\� 6� d� �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ���� ����� � 
�| V ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����8�� )�� �  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    "�j�� , " �
� �  �  
�  m��  ��     ���  �    ]��  ��     ���       h    ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �?�      ��4 �  ��        �&T ���        �        ��        �        ��        �    ��     K�� o��        ��                         ���   	�� ��                                     �                ����             m�����%��   )�8��               18/33 (54%) ek son y   4:52                                                                        2  2     � �
"�'"cV �:c^ �� �� �
 CB �CC �! CI �	C.4 � 
C43 � C5, � C6> �	J�( �J�( � J�8 �J� �J� �J�" � J� |J�$ �k~% � k�5 �c� � � c� � ykj6 qC i C" aC* YC"% aC$" ^c� � ~  c� �!"�$ � ""�6 x#"�$ x$*�3 �%"�3 � &"�E �'�/ �(
�>?)�f � **  +*Lw ,*Rw  -*@  *KWP  *RgX 0*KOP  *Rg � 2*Fw �3*8w � 4*Gw � 5*Pw 6*Fw7*8 8*D_09*
P :*CgX ;*GoX  *KOX  *KOX  *KOP  *Rg                                                                                                                                                                                                                         �� R P               
       �     N P E e  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    �)2�� ��������������������������������������������������������   �4, &  0 9  ���@�@�@��A�	�7��	                                                                                                                                                                                                                                                                                                                          �                                                                                                                                                                                                                                                   B    '     �  D�J    	                                 ������������������������������������������������������                                                                                                                    	                 �      �      �                  �     ~    	  
 	 
 	 	 ���� ����������������� ����������� ����������� ���� ������������������������������� � ����� ���������� �� ��� �� ������ � �������������   �������������� ������������� � ��������������� ����������� �� ��������������������� ��                                $    !    ��  H�J     3�  	                           ������������������������������������������������������                                                                                                                                          �  �     �      �        �    ��              
 	  
	 
 	 	 ����������� �   ����  �������������������������� ���������  ���������� ������� �����   � �� ����� ���������������� ����������� �������� ����  ���������� �������������������� �� ������������������������  ���            x                                                                                                                                                                                                                                                            
                                                 �             


           �   }�         wwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwww , J >               	                  � ��2 �e�                                                                                                                                                                                                                                                                                    �Y  Y              e                  e                  c                                                                                                                                                                                                                                                                                                                                                                                                         � (� �  � (��  � <��  � <��  � (��  JcU  ���������� �����������W�����������������*������                ���� ���        	 	 �   & AG� �  �                 �                                                                                                                                                                                                                                                                                                                                      p B C    �          &             !��                                                                                                                                                                                                                            Y   �� �� ����      �� B 	     ���� ����������������� ����������� ����������� ���� ������������������������������� � ����� ���������� �� ��� �� ������ � �������������   �������������� ������������� � ��������������� ����������� �� ��������������������� ������������� �   ����  �������������������������� ���������  ���������� ������� �����   � �� ����� ���������������� ����������� �������� ����  ���������� �������������������� �� ������������������������  ���             $�������������������˻���������̫�������ʻ������j˻�e���h��fW��jf������̻�j�fUx�f�fffffffffffffff������f�ffgWfff�ffffffffffffffff��������j��̶̻�lV˻fW˫�U��u��˻�������������������������˻��������������������ʺ�˪������������fvf�e�f�fl��jeUfeŘffffffffffffffffffff���i��Vg��ffffffffffffffffffffff�fff�ff�ffhfff�fffffffffe�i�fk��ff�jfffkfffjfffjff�ifffl��������˻������˻�������˪������ʻ�������˺����ʺ���������������fffVf�l�i�x�UʅjYl��Z���WZlvUv�ffff��f�����WxUWwu��Wu���u{fhUZ�ffffU��f��u�uX�[Yu\xwWYwf�W�g�U�ffllfff�fffffffhfffllfffjf�feyXj����������������������������������������������������������������|����ň���uuuXWx�yWy�XuY�xuY�Y�XeUU��UUx�UUW�UUuuUWuu[�u���UyuUUuUUVUUUYuUUUwUUUUUUUUUUUUUUUUUUUgYUke\�j�U�g�UV��UVuyU�u[�kUw[fU�˫�������������������������W������������������������������������W�U�uxW�uw��UX��WY��Wy��U���U���wUux��x�ʪ��yuUX��uYWuUUwuU�wwYUUUUuUUW�UUyuUU�UU[�UW�wW��w�hywxX��vZl�[�j�W���w���XYi�w�j�uuf�X��������������������������������������������������Ȼ��������ǆU�U���W��uX��U[��Uu�fU�kfY�kfVUkƪ��������˸�fhʩfj��fl�jff�ffflḟ���X���������{���h���U��evl�ZfxVl�u�Z���UU�Vl�[fffffffffffffff����̫��Wy�ˇUUXffkUfffhffffffff$�I    4      *      K                       B     � 
 �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$    `d     �f ��     �f �$ ^$ �@      ����� ��   �����    ����` ��   ����` �$ ^$       �                  ,   ���`���� 
"   )+ �Gl ��  �B I ��? �  ��?  �         ��   '���8 e� / �� e� / �$ ^$  �� �� � U ~�c��     	      ���j�������J���� 9� 9"  ��  yf  y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ""   "! " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               ""   "! " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "! ""! " "" """ "!   " ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     �  �  �  ��  �  �  �  ��  �             �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                   ���������������������  ��  ��  ��  �   �    �          �         �                                                                                                                         �   �   �  �  �  �  ���������  �U4"+�B�*�����"/���  ��� �� �  � �     �               ۲  �!  "  �� �� �  ��� ��  �� �                          	ʐ ��� ��� ڝ��ݩ��ݩ��ݩ��ک�̪��̪��̪������̽� ��� ��T �C                �   �   ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                                                 �               �  �  ��  �   �   �                               ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                      �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                       �   �      ��   �  ��  �  �  �         � �������������  �                                                                                                                                         �� v  w � �  �  �  �  
�  ɨ ̊+�˽"˻"�          4   C   C  4  4  3  3   �   �   �   "  "�� ��   �  ��  ��   w   w�  z�  ��� ��� �˰ ̼� �̰ �̰ �˰ ��� ۸� ��@ EHP 5�P E�P H�P X�  X�  H�  E�  ��  ��  ��� (�� "�� �" �"" """ """   �  ��  �  �  �  �   �                      �  ��� ݼ� w��                                      "   "   "                                     �   �  �  �� �  �  �      �   �       ���� �                                                                                                                                                                                       k}z�gg��j�� 
�� 	�� �� �� 
�� �� ��̻�"+��" 4"  4   D   H   H   �  +  ""    ��       ��  �٠ �ڛ ̸� ̻� �̽ �̀ �ɀ ��0 ��C 4�T H�T H�D �T@ �T  �C  �0  ɚ  ��� ��� �" �"  �"�                 �� �� �� {�             �   �� � � ��� � �  ��                                        �   �   �   "   "   "  !�    ��                                                               �               �  �  ��  �   �   �                    �  �˰ ��� �wp ���                                                                                                                                                                                 �  ��� ܽи�؀  � ˚ �̹�̹�˹�˻ܻ��ܘ��܉���D���U�D�J�N T�� D�  T�  �  ��  �� �� ,ث"���"��� ���۝� {�� ��  ��� ��(�������� ˸� ɀ  ��  ��� �̀ �̈ �� ���虎�(���"��� ��� � �/�����              �   �   �   �   �                              � � �  (�  .   .   )�  )�  �   �                 �  ��  �   �  �                      �               �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                                  �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �                   �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                ��� ���� ��                                                                                                                                                                                                  �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �           �  �   �   ��  �            �   �   �   ��                               �� " ��   "             ���� ��� ����                            �    � �  ��                  ���                                                                                                                                                                          �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��                              �                        ���� ��� ����                      �  �� ��  �    � ���                                                                                                                                                                                             	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                                                 �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������             ��  �   ��  �                ���                                                                                                                                                                                             	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��               �� ��������p��}`         �  ��  �  �  ��  �      ��  �              ���  ��                �������  ���    � ��  �   ��  �                    �     �                                                                                                                                                                                                            �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                                                    �   �   �   �   �   �                                                                                                                                                �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(����������������� � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(����������������� 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5���������������� x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x���������������� w w x y�������H���������������������������������H������yxww����������������  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(���������������� , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+���������������� 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5���������������� =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=����������������     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( ���������������� � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � ����������������� � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � ����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
"�'"cV �:c^ �� �� �
 CB �CC �! CI �	C.4 � 
C43 � C5, � C6> �	J�( �J�( � J�8 �J� �J� �J�" � J� |J�$ �k~% � k�5 �c� � � c� � ykj6 qC i C" aC* YC"% aC$" ^c� � ~  c� �!"�$ � ""�6 x#"�$ x$*�3 �%"�3 � &"�E �'�/ �(
�>?)�f � **  +*Lw ,*Rw  -*@  *KWP  *RgX 0*KOP  *Rg � 2*Fw �3*8w � 4*Gw � 5*Pw 6*Fw7*8 8*D_09*
P :*CgX ;*GoX  *KOX  *KOX  *KOP  *Rg3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������� ��=�K�X�X�_��B�G�Q�K� � � � � � � � � � �2�0�.�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.�����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������/�.�7� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� ��!�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y�����������������������9�R�G�_�K�X��<�Z�G�Z�Y�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                