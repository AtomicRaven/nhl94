GST@�                                                            \     �                                               �   �                        ���2���z�	 ʱ��������������z���        �h      #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"      �j* , . ���
��
�"   "D�j��
� " ��
  e                                                                               ����������������������������������       ��    =bo 0Q 4g 11  4              	� 
                     �� � �  �                 En� )         88�����������������������������������������������������������������������������������������������������������������������������oo    og     +      '            ��                     	  7  V  	                  �            :8 �����������������������������������������������������������������������������                                ��  �       �   @  #   �   �                                                                                '     E)n�  �    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�9O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �(���Fl,5E���|@ @#�D��E�C�C#�E���Z3��T0 k� �7��;�2d q51DD"3Q  ��H    ������,���E�l, 7E���|@ @#�D��E�C�C�B���Z3��T0 k� �3��7�2d q51DD"3Q  ��H    ������0���E�p
,$9E���|@ BO#�D��E�C�C�B���Z3��T0 k� �/��3�2d q51DD"3Q  ��H    ������8 ���E�t,(=B���|@ BO#�D��E�?�C�B���Z3��T0 k� �+��/�2d q51DD"3Q  ��H    ������C����E�x,,?B���|@ BO#�D��E�?�S�B���Z3��T0 k� �+��/�2d q51DD"3Q  ��H    ������G����E�|,0AB���|@ BO#�D��E�C�S�B���Z3��T0 k� �'��+�2d q51DD"3Q  �H    ������K���E�|,4CB���|@ BO#�D��E�C�S�B���Z3��T0 k� �+��/�2d q51DD"3Q  ��H    ������S���E��8EB���|@ BO#�D��E�G�S�B��Z3��T0 k� �/��3�2d q51DD"3Q  ��H    ������W���E��<GO/�|?�BO#�D��E�K�S�J@�Z3��T0 k� �3��7�2d q51DD"3Q  ��H    ������_���E��@IO/�|?�BO#�D��E�O�3�J@�Z3��T0 k� �7��;�2d q51DD"3Q  ��H    ������c���E��HKO/�|?�BO#�D��E�O�3�J@�Z3��T0 k� �7��;�2d q51DD"3Q  ��H    ������o���E��POO/�|?�BO#�D��E�W�3�J@#�Z3��T0 k� �;��?�2d q51DD"3Q  ��H    ������s���E��TQO/�|?�BO#�D��E�W�3�E +�Z3��T0 k� �;��?�2d q51DD"3Q  ��H    ������{��w�E��\RO/�|?�BO#�D��E�W�#�E /�Z3��T0 k� �;��?�2d q51DD"3Q  ��H    ��������o�E��`TO/�|?�BO#�D��E�[�#�E 3�Z3��T0 k� �?��C�2d q51DD"3Q  ��H    ���������c�E��hVO/�|?�BO#�D��E�[�#�E 7�Z3��T0 k� �?��C�2d q51DD"3Q  ��H    ���������[�E��lXO/�|?�@#�D��E�[�#�E ;�Z3��T0 k� �?��C�2d q51DD"3Q  �H    �����O���S�E��tZO/�|?�@#�D��E�_�#�E ?�Z3��T0 k� �?��C�2d q51DD"3Q ��O    �����O��C�E����]O/�|?�@#�D��"E�_�#�E G�Z3��T0 k� �;��?�2d q51DD"3Q ��O    �����O��;�E����^O/�|?�@#�D��#E�_�#�E0K�Z3��T0 k� �7��;�2d q51DD"3Q ��O    �����O��3�E����`O/#�|?�@#�D��$E�_�##�E0O�Z3��T0 k� �7��;�2d q51DD"3Q ��O    �����O��'�E����aO/#�|?�BO#�D��%E�_�##�E0S�Z3��T0 k� �3��7�2d q51DD"3Q ��O    �����O���E����cO/'�|?�BO#�D��'E�_�#�E0W�Z3��T0 k� �/��3�2d q51DD"3Q ��O    �����O���E����dO/'�|?�BO#�D��(E�[�'�E0[�Z3��T0 k� �/��3�2d q51DD"3Q ��O    �����O���E��ܨeO/+�|?�BO#�D��)E�[�'�E0[�Z3��T0 k� �+��/�2d q51DD"3Q ��O    �����O���E��ܰfO/+�|?�BO#�D��+E�[�+�E0_�Z3��T0 k� �+��/�2d q51DD"3Q �O    �������� ��E��ܼhO//�|?�BO#�A��-D?W�/�E0d Z3��T0 k� �'��+�2d q51DD"3Q
 �O    ����������CN���iO//�|?�BO#�A��/D?W�/�JphZ3��T0 k� �#��'�2d q51DD"3Q
 ��O   ����������CN� ��jO/3�|?�BO#�A��0D?W�3�JplZ3��T0 k� �#��'�2d q51DD"3Q ��O    ����������CN� ��kE�3�|?�BO#�A��2D?S�3�JplZ3��T0 k� ���#�2d q51DD"3Q ��O    ����������CN���lE�7�|?�BO#�A��3D?S�7�JppZ3��T0 k� ���#�2d q51DD"3Q ��O    ����������CN���mE�7�|?�BO#�A��4D?O�7�JptZ3��T0 k� ����2d q51DD"3Q ��O    ����������CN���mE�;�|?�BO#�A��5D?O�;�Jpx
Z3��T0 k� ����2d q51DD"3Q ��O    ����������CN���nE�?�|?�BO#�A� 7D?K� ;�JpxZ3��T0 k� ����2d q51DD"3Q ��O    ����������CN���nE�?�|?�BO#�A� 8D?K� ?�Jp|Z3��T0 k� ����2d q51DD"3Q ��O    ����������CN�}oE�C�|?�BO#�A�9D?G� ?�Jp�Z3��T0 k� ����2d q51DD"3Q ��O    ����������CN�}oE�C�|?�BO#�A�:D?G� C�Jp�Z3��T0 k� ���2d q51DD"3Q ��O    ����������CN�}pE�G�|?�BO#�A�;D?C� C�Jp�Z3��T0 k� ���2d q51DD"3Q ��O    �����������CN�}pE�G�|?�BO#�A�=DO?� G�Jp�Z3��T0 k� ���2d q51DD"3Q ��O    �����������C^�} pE�K�|?�BO#�A�>DO;� G�Jp�Z3��T0 k� ���2d q51DD"3Q ��O    ����������C^��(pE�K�|?�BO#�A�?DO;� G�Jp�Z3��T0 k� ���2d q51DD"3Q ��O    ���������s�C^��0pE�O�|?�BO#�A�@DO7� K�Jp�Z3��T0 k� ����2d q51DD"3Q ��O    ���������k�C^��8pE�O�|?�BO#�A�ADO3� K�Jp�Z3��T0 k� ����2d q51DD"3Q ��O    ��������c�C^��<pE�S�|?�BO#�A�BDO/� O�Jp�Z3��T0 k� ����2d q51DD"3Q ��O    ��������[�C^��DpE�S�|?�BO#�A�CDO/� O�Jp�Z3��T0 k� �����2d q51DD"3Q ��O    ��������S�C^��LpE�S�|?�BO#�A�DDO+� O�Jp�Z3��T0 k� �����2d q51DD"3Q ��O    ��������K�C^��PoE�W�|?�BO#�A�EDO'� S�Jp�Z3��T0 k� ������2d q51DD"3Q ��O    ��������C�C^��XoE�W�|?�BO#�A�FDO#� P Jp�Z3��T0 k� ������2d q51DD"3Q ��O    ������ �7�C^��`oE�W�|?�BO#�A�GDO� T Jp�Z3��T0 k� ������2d q51DD"3Q ��O    ������ �/�C^��dnE�W�|?�BO#�A�HD_� TJp� Z3��T0 k� ������2d q51DD"3Q ��O    �������'�Cn��lmE�W�|?�BO#�A�ID_� TJp�"Z3��T0 k� ������2d q51DD"3Q ��O    ��������Cn��pmE�W�|?�BO#�A�JD_� XJp�#Z3��T0 k� ������2d q51DD"3Q ��O    ��������Cn��xlE�W�|?�BO#�A�KD_� XJp�$Z3��T0 k� ������2d q51DD"3Q ��O    ��������Cn��|lC�W�|?�BO#�A�LD_� XJp�%Z3��T0 k� ������2d q51DD"3Q ��O    �������Cn���kC�W�|?�BO#�A�ME�� \Jp�&Z3��T0 k� ������2d q51DD"3Q ��O    ������ ��Cn���jC�W�|?�BO#�A�NE�� \Jp�'Z3��T0 k� ������2d q51DD"3Q ��O    �����0 ��Cn���iC�S�|?�BO#�A� OE��� \Jp�(Z3��T0 k� ������2d q51DD"3Q ��O    �����0 ��Cn���hC�S�|?�BO#�A� PE��� `Jp�)Z3��T0 k� ������2d q51DD"3Q ��O    �����?���Cn���gE�S�|?�BO#�A� PE�� `	Jp�*Z3��T0 k� ������2d q51DD"3Q ��O    �����?���Cn�
��fE�O�|?�BO#�A�$QE�� `	Jp�+Z3��T0 k� ������2d q51DD"3Q ��O    �����?���Cn���eE�O�|?�BO#�A�$RE�� d
Jp�,Z3��T0 k� ������2d q51DD"3Q ��O    �����?���E� ��dE�K�|?�BO#�A�$SE�� dJp�-Z3��T0 k� ������2d q51DD"3Q ��O    �����?���E� ��cE�K�|?�BO#�A�$TE�� dJp�.Z3��T0 k� ������2d q51DD"3Q ��O    �����?���E� ��bE�G�|?�BO#�A�(TE�߷ hJp�/Z3��T0 k� ������2d q51DD"3Q ��O    �����?���E�]�aE�G�|?�BO#�A�(UE�۸ hJp�0Z3��T0 k� ������2d q51DD"3Q ��O    �����?���E�]�`E�C�|?�BO#�A�(VE�׸ hJp�1Z3��T0 k� ������2d q51DD"3Q ��O    �����?�/��E� ]�_E�?�|?�BO#�A�(WE�ӹ hJp�2Z3��T0 k� ������2d q51DD"3Q ��O    �����?�/��E��]�^E�?�|?�BO#�A�,XE�Ϻ lJp�3Z3��T0 k� ������2d q51DD"3Q $�O    �����O�/��E��]�^D?;�|?�BO#�A�,Xd�˺ lJp�4Z3��T0 k� ������2d q51DD"3Q ��O    �����O�/��E��]�]D?7�|?�BO#�A�,Yd�ǻ lJp�4Z3��T0 k� ������2d q51DD"3Q ��O    �����O�/��E��]�\D?7�|?�BO#�A�,Zd�ü pJp�5Z3��T0 k� ������2d q51DD"3Q ��O   �����O�/��E��]�[D?3�|?�BO#�A�0Zd��� pJp�6Z3��T0 k� ������2d q51DD"3Q ��O    �����O�/��E��]�ZD?/�|?�BO#�A�0[d��� pJp�7Z3��T0 k� ������2d q51DD"3Q ��O    �����O�/�E��]�YE�+�|?�BO#�A�0\d��� pJp�8Z3��T0 k� ������2d q51DD"3Q ��O    �����O�/{�E��m�XE�'�|?�BO#�A�0\d��� tJp�8Z3��T0 k� ������2d q51DD"3Q ��O    �����O�/w�C��m�XE�#�|?�BO#�A�0]d��� tJp�9Z3��T0 k� ������2d q51DD"3Q ��O    �����O�/o�C��m�WE�#�|?�BO#�A�4^e�� tJp�:Z3��T0 k� ������2d q51DD"3Q ��O    �����O�/k�C��m�VE��|?�BO#�A�4^e�� tJp�;Z3��T0 k� ������2d q51DD"3Q ��O    �����O�/c�C��m�UE��|?�BO#�A�4_e�� xJp�<Z3��T0 k� ������2d q51DD"3Q ��O    �����_�/_�C��m�UE��|?�BO#�A�4`e�� xJp�<Z3��T0 k� ������2d q51DD"3Q ��O    �����_�/[�C��m�TE��|?�BO#�A�4`e�� xJp�=Z3��T0 k� ������2d q51DD"3Q ��O    �����_�/S�C��n SE��|?�BO#�A�8ae�� xJp�>Z3��T0 k� ������2d q51DD"3Q ��O    �����_� /O�C��nRE��|?�BO#�A�8ae�� xJp�>Z3��T0 k� ������2d q51DD"3Q ��O    �����_� /K�C��nRF�|?�BO#�A�8bF�� |Jp�?Z3��T0 k� ������2d q51DD"3Q ��O    �����_��/C�C��nQF�|?�BO#�A�8bF�� |Jp�@Z3��T0 k� ������2d q51DD"3Q ��O    �����_��/C�C��nPF�|?�BO#�A�8cF�� |Jp�@Z3��T0 k� ������2d q51DD"3Q ��O    �����_��/?�C��nPF�|?�BO#�A�<dF�� |Jp�AZ3��T0 k� �����2d q51DD"3Q $�O    �����_��/?�C��nOF��|?�BO#�A�<dF�� |Jp�BZ3��T0 k� �����2d q51DD"3Q ��O   �����_��/?�d~��nNF��|?�BO#�A�<eF�� �Jp�BZ3��T0 k� �����2d q51DD"3Q ��O    �����_��/;�d~��nNF��|?�BO#�A�<eE��� �Jp�CZ3��T0 k� �����2d q51DD"3Q ��O    �����o��/;�d~��n ME���|?�BO#�A�<fE��� �Jp�DZ3��T0 k� �����2d q51DD"3Q ��O   �����o��/7�d~��n$LE���|?�BO#�A�<fE��� �Jp�DZ3��T0 k� ������2d q51DD"3Q ��O    �����o��/7�d~��n(LE���|?�BO#�A�@gE��� �Jp�EZ3��T0 k� ������2d q51DD"3Q ��O    �����o��/7�d~��n,KE���|?�BO#�A�@gE��� �Jp�EZ3��T0 k� ������2d q51DD"3Q ��O    �����o{�/3�d~��n,KE���|?�BO#�A�@hE��� �Jp�FZ3��T0 k� ������2d q51DD"3Q
 $�O    �����ow�/3�d���n0JE���|?�BO#�A�@hE��� �Jp�GZ3��T0 k� ������2d q51DD"3Q
 ��O    �����oo�/3�d���n4JE���|?�BO#�A�@iE��� �Jp�GZ3��T0 k� ������2d q51DD"3Q
 ��O    �����ok�/3�d���n8IE���|?�BO#�A�@iE��� �Jp�HZ3��T0 k� ������2d q51DD"3Q
 ��O    �����oc�/3�d���n8HE���|?�BO#�A�DjE��� �Jp�HZ3��T0 k� ������2d q51DD"3Q
 ��O    �����o_�/3�d���n<HE���|?�BO#�A�DjE��� �Jp�IZ3��T0 k� ������2d q51DD"3Q
 ��O    �����oW�/3�d���n@GB���|?�BO#�A�DjE��� � Jp�IZ3��T0 k� ������2d q51DD"3Q
 ��O    �����?S�/3�d���n@GB���|?�BO#�A�DkE��� � Jp�JZ3��T0 k� ������2d q51DD"3Q
 ��O    �����?K�/3�C���nDFB���!�?�BO#�A�DkE��� �!Jp�Jb���T0 k� ������2d q51DD"3Q	 ��O    �����?G�/3�C���nHFB���!�?�BO#�A�DlE��� �!Jp�Kb���T0 k� ������2d q51DD"3Q	 ��O    �����??�/3�C���nHEB���!�?�BO#�A�DlB��� �!Jp�Kb���T0 k� ������2d q51DD"3Q	 ��O   �����?7�/3�C���nLEB���!�?�BO#�A�HmB��� �"Jp�Lb���T0 k� ������2d q51DD"3Q	 ��O    �����?3�/3�C���nPDB���!�?�BO#�A�HmB��� �"Jp�Lb���T0 k� �����2d q51DD"3Q ��O    �����?+�3�C���nPDB���!�?�BO#�A�HmB��� �"Jp�Mb���T0 k� �����2d q51DD"3Q ��O    �����?'�3�C���nTCB���!�?�BO#�A�HnB��� �#Jp�Mb���T0 k� �����2d q51DD"3Q ��O    �������3�C���nXCB���!�?�BO#�A�HnB��� �#Jp�Nb���T0 k� �����2d q51DD"3Q ��O    �������7�C���nXBB���!�?�BO#�A�Hn@�� �$Jq Nb���T0 k� �����2d q51DD"3Q ��O    �������7�E>��n\BB���!�?�BO#�A�Ho@�� �$Jq Ob���T0 k� �����2d q51DD"3Q ��O    �������7�E>��n\BB��!�?�BO#�A�Ho@�� �$Jq Ob���T0 k� �����2d q51DD"3Q ��O    �������_7�E>��n`AB��|?�BO#�A�Lp@�� �$Jq OZ3��T0 k� �����2d q51DD"3Q ��O    ��������_7�E>��ndAB��|?�BO#�A�Lp@�� �%Jq PZ3��T0 k� �����2d q51DD"3Q ��O    ��������_7�E>��^d@B��|?�BO#�A�LpB��� �%JqPZ3��T0 k� �����2d q51DD"3Q ��O    ��������_7�E>��^h@B��|?�BO#�A�LqB��� �%JqQZ3��T0 k� ������2d q51DD"3Q ��O    ��������_7�E>��^h?E��|?�BO#�A�LqB��� �&JqQZ3��T0 k� ������2d q51DD"3Q �O    ��������?7�S���^l?E��|?�BO#�A�LqB��� �&JqQZ3��T0 k� ������2d q51DD"3Q ��O    ��������?7�S���^l?E��|?�BO#�A�LrB��� �&JqRZ3��T0 k� ������2d q51DD"3Q ��O    ��������?;�S���^p>E��|?�BO#�A�LrO�� �'JqRZ3��T0 k� ������2d q51DD"3Q ��O    ��������?;�S����p>E��|?�BO#�A�LrO�� �'JqSZ3��T0 k� ������2d q51DD"3Q  ��O   ��������?;�S����t=L�|?�BO#�A�PsO�� �'JqSZ3��T0 k� ������2d q51DD"3Q  ��O    �����n��?;�S����t=L�|?�BO#�A�PsO�� �'JqSZ3��T0 k� ������2d q51DD"3Q  ,�O   �����n��?;�S����x<L�!�?�BO#�A�PsO�� �(JqTbs��T0 k� ������2d q51DD"3Q  ��O   �����n��?7�S����x;L�!�?�BO#�A�PtO�� �(JqTbs��T0 k� ������2d q51DD"3Q  ��O    �����n��?7�S����|;L�!�?�BO#�A�PtO�� �(JqTbs��T0 k� ������2d q51DD"3Q  ��O    �����n��?7�S����|:L�!�?�BO#�A�PtO�� �)JqUbs��T0 k� ������2d q51DD"3Q ��O    �����n��?7�S�����9L#�!�?�BO#�A�PtO�� �)JqUbs��T0 k� ������2d q51DD"3Q ��O    �����n��O7�S�����8L#�!�?�BO#�A�PuO�� �)JqUbs��T0 k� ������2d q51DD"3Q ��O    �����n��O7�S�����7L'�!�?�BO#�A�PuO�� �)JqVbs��T0 k� ������2d q51DD"3Q ��O    �����>��O7�S�����6L'�!�?�BO#�A�PuO�� �*JqVbs��T0 k� �����2d q51DD"3Q ��O    �����>��O7�S�����5L+�!�?�BO#�A�TuO�� �*JqVbs��T0 k� �����2d q51DD"3Q ��O    �����>��O7�S�����4L+�!�?�BO#�A�TvO�� �*JqWbs��T0 k� �����2d q51DD"3Q ��O    �����>��O7�S�����3L/�!�?�BO#�A�TvO�� �*JqWbs��T0 k� �����2d q51DD"3Q ��O    �����>��O7�S�����2L�/�|?�BO#�A�TvO�� �*JqWZ3��T0 k� �����2d q51DD"3Q ��O    �����>��O7�S�����0L�/�|?�BO#�A�TwO�� �+JqXZ3��T0 k� �����2d q51DD"3Q ��O    �����>��O7�S�����/L�3�|?�BO#�A�TwO�� �+JqXZ3��T0 k� �����2d q51DD"3Q ��O    �����>��O7�S�����.L�3�|?�BO#�A�TwO�� �+JqXZ3��T0 k� �����2d q51DD"3Q ��O    �����>��O7�S�����,L�3�|?�BO#�A�TwO�� �+JqYZ3��T0 k� �����2d q51DD"3Q ��O    �����>��_7�S�����+L�7�|?�BO#�A�TxO�� �,JqYZ3��T0 k� �����2d q51DD"3Q ��O    �����>��_7�S�����)L�7�|?�BO#�A�TxO�� �,JqYZ3��T0 k� ������2d q51DD"3Q ��O    �����>��_7�S�����(L�;�|?�BO#�A�TxO�� �,JqYZ3��T0 k� ������2d q51DD"3Q ��O    �����>��_3�S�����&L�;�|?�BO#�A�TxO�� �,JqZZ3��T0 k� ������2d q51DD"3Q ��O    �����>��_3�S�����%L�;�|?�BO#�A�XxB��� �,JqZZ3��T0 k� ������2d q51DD"3Q ��O    �����>��_3�S�����#L�?�|?�BO#�A�XyB��� �-JqZZ3��T0 k� ������2d q51DD"3Q ��O    �����>��_3�S�����!L�?�|?�BO#�A�XyB��� �-JqZZ3��T0 k� ������2d q51DD"3Q ��O    �����>��_3�S����� L�?�|?�BO#�A�XyB��� �-Jq[Z3��T0 k� ������2d q51DD"3Q ��O    �����>��_/�S�����L�C�|?�BO#�A�XyB��� �-Jq[Z3��T0 k� ������2d q51DD"3Q  ��O    �����>��_/�S�����L�C�|?�BO#�A�Xz@�� �-Jq[Z3��T0 k� ������2d q51DD"3Q  ��O    �����>��_/�S�����L�C�|?�BO#�A�Xy@�� �.Jq[Z3��T0 k� ������2d q51DD"3Q  ��O    �����>��o+�S�����L�G�|?�BO#�A�Xy@�� �.Jq\Z3��T0 k� ������2d q51DD"3Q  ��O    �����>��o+�S�����L�G�|?�BO#�A�Xy@�� �.Jq\Z3��T0 k� ������2d q51DD"3Q  /�O    �����>��o+�S�����L�G�|?�BO#�A�Xy@�� �.Jq\Z3��T0 k� ������2d q51DD"3Q  ��O    �����>��o'�S�����L�G�|?�BO#�A�Xx@�� �.Jq\Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��o'�S�����L�K�|?�BO#�A�Xx@�� �.Jq]Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��o#�S�����L�K�|?�BO#�A�Xx@�� �/Jq]Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��o#�S�����L�K�|?�BO#�A�Xx@�� �/Jq]Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��o�S�����
L�O�|?�BO#�A�\w@�� �/Jq]Z3��T0 k� ������2d q51DD"3Q  ��O   �����N��o�S�����L�O�|?�BO#�A�\w@�� �/Jq^Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��o�S�����L�O�|?�BO#�A�\w@�� �/Jq ^Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��o�S�����L�O�|?�BO#�A�\w@�� �/Jq ^Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��o�S�����L�S�|?�BO#�A�\v@�� �0Jq ^Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��_�S������L�S�|?�BO#�A�\v@�� �0Jq ^Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��_�S������L�S�|?�BO#�A�\v@�� �0Jq _Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��_�S������L�S�|?�BO#�A�\v@�� �0Jq _Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��_�S������L�W�|?�BO#�A�\v@�� �0Jq _Z3��T0 k� ������2d q51DD"3Q  ��O    �����N��^��S������L�W�|?�BO#�A�\u@�� �0Jq _Z3��T0 k� ������2d q51DD"3Q  ��O    �����N�����S������L�W�|?�BO#�A�\u@�� �0Jq _Z3��T0 k� ������2d q51DD"3Q  ��O    �����N�����S������L�W�|?�BO#�A�\u@�� �1Jq _Z3��T0 k� ������2d q51DD"3Q  ��O    �����N����S���~��L�[�|?�BO#�A�\u@�� �1Jq$`Z3��T0 k� ������2d q51DD"3Q  ��O    �����N����S���~��L�[�|?�BO#�A�\u@�� �1Jq$`Z3��T0 k� ������2d q51DD"3Q  ��O    �����N����S���~��L�[�|?�BO#�A�\t@�� �1Jq$`Z3��T0 k� ������2d q51DD"3Q  ��O    �����N����S���~��L�_�|?�BO#�A�\t@�� �1Jq$`Z3��T0 k� ������2d q51DD"3Q  ��O    �����N����S���~��L�_�|?�BO#�A�`t@�� �1Jq$aZ3��T0 k� ������2d q51DD"3Q  ��O    �����N���߮S���~��L_�|?�BO#�A�`t@�� �2Jq$aZ3��T0 k� ������2d q51DD"3Q  ��O    �����N���߭S���~��L_�|?�BO#�A�`t@�� �2Jq$aZ3��T0 k� ������2d q51DD"3Q  ��O    �����N���߭S���~��L_�|?�BO#�A�`t@�� �2Jq$aZ3��T0 k� ������2d q51DD"3Q  ��O    �����N���۬S���~��Lc�|?�BO#�A�`s@�� �2Jq$aZ3��T0 k� ������2d q51DD"3Q  ��O    �����N���۬S���~��Lc�|?�BO#�A�`s@�� �2Jq$aZ3��T0 k� ������2d q51DD"3Q  ��O    �����N���׫S���n��Lc�|?�BO#�A�`s@�� �2Jq(bZ3��T0 k� ������2d q51DD"3Q  ��O    �����N���ӪS���n��BOc�|?�BO#�A�`s@�� �2Jq(bZ3��T0 k� ������2d q51DD"3Q  ��O    �����N���ӪS���n��BOc�|?�BO#�A�`s@�� �2Jq(bZ3��T0 k� ������2d q51DD"3Q  ��O    �����N���өS���n��BOg�|?�BO#�A�`s@�� �2Jq(bZ3��T0 k� ������2d q51DD"3Q  ��O   �����N۾^ϩS���n��BOg�|?�BO#�A�`r@�� �3Jq(bZ3��T0 k� ������2d q51DD"3Q  ��O    �����N۽^˨S���n��BOg�|?�BO#�A�`r@�� �3Jq(bZ3��T0 k� ������2d q51DD"3Q  ��O    �����Nۼ^ǧS���n��BOg�|?�BO#�A�`r@�� �3Jq(bZ3��T0 k� ������2d q51DD"3Q  ��O    �����Nۻ^ǧS���n��BOg�|?�BO#�A�`r@�� �3Jq(cZ3��T0 k� ������2d q51DD"3Q  ��O    �����Nۺ^æS���n��BOk�|?�BO#�A�`r@�� �3Jq(cZ3��T0 k� ������2d q51DD"3Q  ��O    �����N۹NæS���n��BOk�|?�BO#�A�`r@�� �3Jq(cZ3��T0 k� ������2d q51DD"3Q  ��O    �����N۸N��S���^��BOk�|?�BO#�A�`r@�� �3Jq(cZ3��T0 k� ������2d q51DD"3Q  ��O    �����N۷N��S���^��BOk�|?�BO#�A�`r@�� �3Jq(cZ3��T0 k� ������2d q51DD"3Q  ��O    �����N۶N��S���^��BOk�|?�BO#�A�`q@�� �3Jq(cZ3��T0 k� ������2d q51DD"3Q  ��O    �����N۵N��S���^��BOk�|?�BO#�A�`q@� �4Jq(cZ3��T0 k� ������2d q51DD"3Q  ��O    �����Nߴ���S��^��BOo�|?�BO#�A�`q@� �4Jq,cZ3��T0 k� ������2d q51DD"3Q  ��O    �����>߳���S�{���BOo�|?�BO#�A�`q@� �4Jq,dZ3��T0 k� ������2d q51DD"3Q  ��O    �����>߲���S�{���BOo�|?�BO#�A�dq@{� �4Jq,dZ3��T0 k� ������2d q51DD"3Q  ��O    �����>߱���S�w���BOo�|?�BO#�A�dq@{� �4Jq,dZ3��T0 k� ������2d q51DD"3Q  ��O    �����>߰���S�w���BOo�|?�BO#�A�dq@w� �4Jq,dZ3��T0 k� ������2d q51DD"3Q  ��O   �����>߯���S�s���BOo�|?�BO#�A�dq@w� �4Jq,dZ3��T0 k� ������2d q51DD"3Q  ��O    �����>߮���S�s���BOo�|?�BO#�A�dp@s� �4Jq,dZ3��T0 k� �� �� 2d q51DD"3Q  ��O    �����>߭���S�o�BOs�|?�BO#�A�dp@s� �4Jq,dZ3��T0 k� �� �� 2d q51DD"3Q  ��O    �����>߬���S�o�BOs�|?�BO#�A�dp@s� �4Jq,dZ3��T0 k� �� �� 2d q51DD"3Q  ��O    �����>߫���S�k�>��BOs�|?�BO#�A�dp@o� �4Jq,eZ3��T0 k� ����2d q51DD"3Q  ��O    �����>ߪ���S�k�>��BOs�|?�BO#�A�dp@o� �5Jq,eZ3��T0 k� ����2d q51DD"3Q  ��O    �����>ߩ���S�g�>��BOs�|?�BO#�A�dp@o� �5Jq,eZ3��T0 k� ����2d q51DD"3Q  ��O   �����nߨ���S�g�>��BOs�|?�BO#�A�dp@k� �5Jq,eZ3��T0 k� ����2d q51DD"3Q  ��O    �����nۧ���S�g�>��BOs�|?�BO#�A�dp@k� �5Jq,eZ3��T0 k� ����2d q51DD"3Q  ��O    �����nۦ���S�c�	���BOw�|?�BO#�A�dp@g� �5Jq,eZ3��T0 k� ����2d q51DD"3Q  ��O    �����nۥ���S�c�	���BOw�|?�BO#�A�dp@g� �5Jq,eZ3��T0 k� ����2d q51DD"3Q  ��O    �����nפ���S�_�	���BOw�|?�BO#�A�do@g� �5Jq,eZ3��T0 k� ����2d q51DD"3Q  ��O    �����nף���S�_�	���BOw�|?�BO#�A�do@c� �5Jq0eZ3��T0 k� ����2d q51DD"3Q  ��O    �����nס���S�[�	���BOw�|?�BO#�A�do@c� �5Jq0eZ3��T0 k� ����2d q51DD"3Q  ��O    �����^ס���S�[�	Λ�BOw�|?�BO#�A�do@_� �5Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^נ���S�[�	Λ�BOw�|?�BO#�A�do@_� �5Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^ӟ���S�W�	Λ�BOw�|?�BO#�A�do@[� �5Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^Ӟ���S�W�	Λ�BO{�|?�BO#�A�do@[� �5Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^ϝ���S�S�	Λ�BO{�|?�BO#�A�do@W� �6Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^ϛ��S�S�>��BO{�|?�BO#�A�do@W� �6Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^˚��S�S�>��BO{�|?�BO#�A�do@W� �6Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O   �����^Ǚ��S�O�>��BO{�|?�BO#�A�do@S� �6Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^Ø��S�O�>��BO{�|?�BO#�A�dn@S� �6Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^����S�O�>��BO{�|?�BO#�A�dn@O� �6Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^����S�K�>��BO{�|?�BO#�A�dn@O� �6Jq0fZ3��T0 k� ����2d q51DD"3Q  ��O    �����^���S�K�>��BO{�|?�BO#�A�dn@O� �6Jq0gZ3��T0 k� ����2d q51DD"3Q  ��O    �����^���S�K�>��BO�|?�BO#�A�dn@K� �6Jq0gZ3��T0 k� ����2d q51DD"3Q  ��O   �����N��{�S�G�>��BO�|?�BO#�A�dn@K� �6Jq0gZ3��T0 k� ����2d q51DD"3Q  ��O    �����N��{�S�G�>��BO�|?�BO#�A�hn@G� �6Jq0gZ3��T0 k� ����2d q51DD"3Q  ��O    �����N��w�S�G�>��BO�|?�BO#�A�hn@G� �6Jq0gZ3��T0 k� ����2d q51DD"3Q  ��O    �����N��w�S�C�>��BO�|?�BO#�A�hn@G� �6Jq0gZ3��T0 k� ����2d q51DD"3Q  ��O    �����N��w�S�C�N��BO�|?�BO#�A�hn@C� �6Jq0gZ3��T0 k� ����2d q51DD"3Q  ��O    �����N��s�S�C�N��BO�|?�BO#�A�hn@C� �6Jq0gZ3��T0 k� ��	��	2d q51DD"3Q  ��O    ��������s�S�?�N��BO�|?�BO#�A�hn@C� �6Jq0gZ3��T0 k� ��	��	2d q51DD"3Q  ��O    ��������o�S�?�N��BO�|?�BO#�A�hn@?� �6Jq4gZ3��T0 k� ��	��	2d q51DD"3Q  ��O    ��������o�S�?�N��BO�|?�BO#�A�hn@?� �7Jq4gZ3��T0 k� ��	��	2d q51DD"3Q  ��O    ��������o�S�?�N��BO�|?�BO#�A�hn@?� �7Jq4gZ3��T0 k� ��
��
2d q51DD"3Q  ��O    ��������k�S�;�N��BO��|?�BO#�A�hm@;� �7Jq4gZ3��T0 k� ��
��
2d q51DD"3Q  ��O    ��������k�S�;�N��BO��|?�BO#�A�hm@;� �7Jq4hZ3��T0 k� ��
��
2d q51DD"3Q  ��O    ��������k�S�;�N��BO��|?�BO#�A�hm@;� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    �������g�S�7�N��BO��|?�BO#�A�hm@7� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    ������{�g�S�7�N��BO��|?�BO#�A�hm@7� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    ������w�c�S�7�N��BO��|?�BO#�A�hm@7� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    ������s�c�U>7�N��BO��|?�BO#�A�hm@7� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    ������o�c�U>3�N��BO��|?�BO#�A�hm@3� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    ������o�_�U>3�N��BO��|?�BO#�A�hm@3� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    ������k�_�U>3�N��BO��|?�BO#�A�hm@3� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    �����g�_�U>3�N��BO��|?�BO#�A�hm@/� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    �����c�[�U>/�N��BO��|?�BO#�A�hm@/� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    �����_�[�U>/�N��BO��|?�BO#�A�hm@/� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O   �����[�[�U>/�N��BO��|?�BO#�A�hm@/� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    �����[�[�U>/�N��BO��|?�BO#�A�hm@+� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    �����W�W�CN/�N��BO��|?�BO#�A�hm@+� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    �����S�W�CN+�N��L��|?�BO#�A�hm@+� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O   �����O�W�CN+�N��L��|?�BO#�A�hm@+� �7Jq4hZ3��T0 k� ����2d q51DD"3Q  ��O    �����O�W�CN+�N��L��|?�BO#�A�hm@'� �8Jq4iZ3��T0 k� ����2d q51DD"3Q  ��O    �����K�W�CN+�N��L��|?�BO#�A�hm@'� �8Jq4iZ3��T0 k� ����2d q51DD"3Q  ��O    �����G�W�E>'�N��L��|?�BO#�A�hl@'� �8Jq4iZ3��T0 k� ����2d q51DD"3Q  ��O    �����C�W�E>'�N��L��|?�BO#�A�hl@'� �8Jq4iZ3��T0 k� ����2d q51DD"3Q  ��O    �����C�S�E>'�N��L��|?�BO#�A�hl@#� �8Jq4iZ3��T0 k� ����2d q51DD"3Q  ��O    �����?��S�E>'�N��L��|?�BO#�A�hl@#� �8Jq4iZ3��T0 k� ����2d q51DD"3Q  ��O    �����;��S�E>'�N��L��|?�BO#�A�hl@#� �8Jq4iZ3��T0 k� ����2d q51DD"3Q  ��O    �����;��S�E.'�N��L��|?�BO#�A�hl@#� �8Jq4iZ3��T0 k� ����2d q51DD"3Q  ��O    �����7��O�E.'�N��L��|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    �����3��O�E.'�N��L��|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    �����3��O�E.'�N��L��|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    �����/��O�E.'�N��L��|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    �����+�O�B�'�N��L���|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    �����+�O�B�'�N��L���|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    �����'�O�B�'�N��L���|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    �����'�O�B�'�N��L���|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    �����#�O�B�+�N��L���|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    ������ �K�E.+�>��L���|?�BO#�A�hl@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    ������ �K�E.+�>��L���|?�BO#�A�ll@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    ������ �K�E./�>��L���|?�BO#�A�ll@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    ������ �K�E./�>��L���|?�BO#�A�ll@� �8Jq8iZ3��T0 k� ����2d q51DD"3Q  ��O    ������ �K�E./�>��L���|?�BO#�A�ll@� �8Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    ������ nK�E3�>��L���|?�BO#�A�ll@� �8Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    ������ nK�E7�>��L���|?�BO#�A�ll@� �8Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    ������ nK�E7�>��L���|?�BO#�A�ll@� �8Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    ������ nK�E;�>��L���|?�BO#�A�ll@� �8Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    ������ nK�E;�>��L���|?�BO#�A�ll@� �8Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������K�B�?�>��L���|?�BO#�A�ll@� �8Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������K�B�?����L���|?�BO#�A�ll@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������K�B�C����L���|?�BO#�A�ll@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������K�B�C����L���|?�BO#�A�ll@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������K�B�C����L���|?�BO#�A�ll@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    ������ nK�K�G����L���|?�BO#�A�ll@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������� nK�K�G����L���|?�BO#�A�ll@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������� nK�K�K����L���|?�BO#�A�lk@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������� nK�K�K����L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������� nK�K�K�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������� �K�K�O�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �������� �K�K�O�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����M�� �K�K�S�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����M� �K�K�S�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����M� �K�K�S�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����M� �K�K�W�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����M� �K�K�W�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����=� �K�K�W�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����=� �K�K�[�^��L���|?�BO#�A�lk@�� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����=� �K�K�[�^��L���|?�BO#�A�lk@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����=� �K�K�_�^��L���|?�BO#�A�lk@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����=� �K�K�_���L���|?�BO#�A�lk@� �9Jq8jZ3��T0 k� ����2d q51DD"3Q  ��O    �����=� �K�K�_���L���|?�BO#�A�lk@� �9Jq8kZ3��T0 k� ����2d q51DD"3Q  ��O    �����=ߌ �K�K�_���L���|?�BO#�A�lk@� �9Jq8kZ3��T0 k� ����2d q51DD"3Q  ��O    �����=ߍ �K�K�c���L���|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O    �����=ߍ �K�K�c���L���|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O    �����-ߍ �K�K�c���L��|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O    �����-ߍ �K�K�g���L��|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O    �����-ߍ �K�K�g���L��|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O    �����-ێ �K�K�g���L��|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O    �����-ێ �K�K�g���L��|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O   �����-׏ �K�K�g���L��|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O    �����׏ �K�K�g���BO��|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O    �����א �K�K�g���BO��|?�BO#�A�lk@� �9Jq<kZ3��T0 k� ����2d q51DD"3Q  ��O    �����א �K�K�g���BO��!�?�BO#�A�lk@� �9Jq<kbs��T0 k� ����2d q51DD"3Q  ��O    �����ב �K�K�g���BO��!�?�BO#�A�lk@� �9Jq<kbs��T0 k� ����2d q51DD"3Q  ��O    �����ב �K�K�k���BO��!�?�BO#�A�lk@� �9Jq<kbs��T0 k� ����2d q51DD"3Q  ��O    �����ב �K�K�k���BO��!�?�BO#�A�lk@� �9Jq<kbs��T0 k� �� �� 2d q51DD"3Q  ��O    �����ב �K�K�k���BO��!�?�BO#�A�lk@� �9Jq<kbs��T0 k� �� �� 2d q51DD"3Q  ��O    �����ב �K�K�k���BO��!�?�BO#�A�lk@� �9Jq<kbs��T0 k� �� �� 2d q51DD"3Q  ��O    �����ג �K�K�k���L��!�?�BO#�A�lk@� �:Jq<kbs��T0 k� �� �� 2d q51DD"3Q  ��O    �����ے �K�K�k���L��!�?�BO#�A�lk@� �:Jq<kbs��T0 k� ��!��!2d q51DD"3Q  ��O    ������ے �K�K�k���L��!�?�BO#�A�lk@� �:Jq<kbs��T0 k� ��!��!2d q51DD"3Q  ��O    ������ے �K�K�k���L��!�?�BO#�A�lk@� �:Jq<kbs��T0 k� ��!��!2d q51DD"3Q  ��O    ������ߒ �K�K�k���L��!�?�BO#�A�lk@� �:Jq<kbs��T0 k� ��!��!2d q51DD"3Q  ��O    ������ߒ �K�K�k� ���L��|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��"��"2d q51DD"3Q  ��O    ������� �K�K�k� ���L��|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��"��"2d q51DD"3Q  ��O    ������� �K�K�k� ���L��|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��"��"2d q51DD"3Q  ��O    ������� �K�K�k� ���L��|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��"��"2d q51DD"3Q  ��O    ������� �K�K�k� ���L��|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��#��#2d q51DD"3Q  ��O    ������� �K�K�k� ���L��|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��#��#2d q51DD"3Q  ��O    ������� �K�K�k� ���L��|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��#��#2d q51DD"3Q  ��O    ������� �K�K�k� ���L��|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��#��#2d q51DD"3Q  ��O    ������� �K�K�k� ���L��|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��$��$2d q51DD"3Q  ��O    ������� �K�K�k� ���L���|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��$��$2d q51DD"3Q  ��O    ������� �K�K�k� ���L���|?�BO#�A�lk@� �:Jq<kZ3��T0 k� ��$��$2d q51DD"3Q  ��O    �������� �K�K�k� ���L���!�?�BO#�A�lk@� �:Jq<kb���T0 k� ��$��$2d q51DD"3Q  ��O    �������� �K�K�k� ���L���!�?�BO#�A�lk@� �:Jq<kb���T0 k� ��$��$2d q51DD"3Q  ��O    �������� �K�K�k� ���L���!�?�BO#�A�lk@� �:Jq<kb���T0 k� ��%��%2d q51DD"3Q  ��O    ������� �K�K�k� ���L���!�?�BO#�A�lk@� �:Jq<kb���T0 k� ��%��%2d q51DD"3Q  ��O    ������ �K�K�k� ���L���!�?�BO#�A�lk@� �:Jq<kb���T0 k� ��%��%2d q51DD"3Q  ��O    ������ �K�K�k� ���L���!�?�BO#�A�lk@� �:Jq<kb���T0 k� ��%��%2d q51DD"3Q  ��O    ������ �O�K�k� ���L���!�?�BO#�A�lk@� �:Jq<kb���T0 k� ��&��&2d q51DD"3Q  ��O    ������ �O�K�k� ���L���!�?�BO#�A�lk@� �:Jq<lb���T0 k� ��&��&2d q51DD"3Q  ��O    ������ �S�@k� ���L���!�?�BO#�A�lk@� �:Jq<lb���T0 k� ��&��&2d q51DD"3Q  ��O    ������ �S�@k� ���L���!�?�BO#�A�lk@� �:Jq<lb���T0 k� ��&��&2d q51DD"3Q  ��O    ������ �W�@k� ���L���!�?�BO#�A�lk@� �:Jq<lb���T0 k� ��'��'2d q51DD"3Q  ��O    ������� �W�@k� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��'��'2d q51DD"3Q  ��O    ������� �[�@k� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��'��'2d q51DD"3Q  ��O    ������� �[�@k� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��'��'2d q51DD"3Q  ��O    ������� �[�@k� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��(��(2d q51DD"3Q  ��O    ������� �_�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��(��(2d q51DD"3Q  ��O    ������� �_�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��(��(2d q51DD"3Q  ��O    ������� �_�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��(��(2d q51DD"3Q  ��O    ������� �_�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��)��)2d q51DD"3Q  ��O    ������� �_�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��)��)2d q51DD"3Q  ��O    ������� �_�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��)��)2d q51DD"3Q  ��O    ������� �c�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��)��)2d q51DD"3Q  ��O    ������� �c�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��*��*2d q51DD"3Q  ��O    ������� �c�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��*��*2d q51DD"3Q  ��O    ��������c�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��*��*2d q51DD"3Q  ��O    ��������c�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��*��*2d q51DD"3Q  ��O    ��������c�BNk� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��+��+2d q51DD"3Q  ��O    ������#��c�A�k� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��+��+2d q51DD"3Q  ��O    ������#��c�A�k� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��+��+2d q51DD"3Q  ��O    ������#��c�A�k� ���L���|?�BO#�A�lk@� �:Jq<lZ3��T0 k� ��+��+2d q51DD"3Q  ��O    ������v��E��M#E�#��3�E.��C_8}E��6
�7�E�ψZ3��T0 k� �Ö�ǖ2d q51DD"3Q  ��J    ����}�v�{�E��M"E�'��3�E.��C_8}E��7
�;�E�ψZ3��T0 k� �˘�Ϙ2d q51DD"3Q  ��J    ����}|u�{�E���M"E�'��3�E.��C_4}E��7
�;�E�ωZ3��T0 k� �ϙ�ә2d q51DD"3Q  ��J    ����}xt�{�E���M "E�'��3�E.��C_4}E��8
�;�E�ӉZ3��T0 k� �ӛ�כ2d q51DD"3Q  ��J    ����~tt�{�E}��L�!E�+��3�E.��C_4|B��8
�;�E�ӈZ3��T0 k� �ۛ�ߛ2d q51DD"3Q  ��J    ����ts�{�E}����!E�+��3�E.��C_4|B��8
�;�F׈Z3��T0 k� ����2d q51DD"3Q  ��J    �����lr�{�E}���� E�/��3�E��C_0{B��9
�;�FۈZ3��T0 k� �����2d q51DD"3Q  ��J    �����hq�{�E}����E~3��3�E��C_0{B��9
�;�FۈZ3��T0 k� ������2d q51DD"3Q  ��J    �����dq�{�D�����E~3��3�E��C_,zB��:
�;�F߉Z3��T0 k� �����2d q51DD"3Q  ��J    �����`p�{�D�����E~7��3�E��C_,zB��:
�;�E~߉Z3��T0 k� ������2d q51DD"3Q  ��J    �����\o�{�D����E~7��3�E��Co,zE� :
�;�E~�Z3��T0 k� ������2d q51DD"3Q  ��J    �����Xn�{�D����E~;��3�E���Co(yE� :
�;�E~�Z3��T0 k� ������2d q51DD"3Q  ��J    �����Xn�{�D����D�;��3�E���Co$yE�:
�;�E~�Z3��T0 k� ������2d q51DD"3Q  ��J    �����Tm�{�D����D�?��3�E���Co$xE�:
�;�E~�Z3��T0 k� ������2d q51DD"3Q  ��J    �����Lk�{�D����D�C��3�E���CowE�:
�;�E~�Z3��T0 k� ������2d q51DD"3Q  ��J    �����Hj�{�D����D�C��3�E���CovE�:
�;�B�Z3��T0 k� �����2d q51DD"3Q  ��J    �����	�Hj�{�D����D~C��3�E���CovE�:
�;�B�Z3��T0 k� ����2d q51DD"3Q  ��J    �����	�Di�{�D���tD~G��3�E>��CouE�:
�;�B�Z3��T0 k� ����2d q51DD"3Q  ��J    �����	�@h�{�D���lD~G��3�E>��CotE�9
�;�B�Z3��T0 k� ����2d q51DD"3Q  ��J    �����	�@h�{�D���hD~G��3�E>��CosE�9
�;�B�Z3��T0 k� ����2d q51DD"3Q  ��J    �����	�<g�{�D���`D~G��3�E>��CsCO9
�;�F��Z3��T0 k� �����2d q51DD"3Q  ��J    �����	�8f�{�D���XN�G��3�E>��CsCO8
�;�F��Z3��T0 k� ����2d q51DD"3Q  �J    �����	�4e�{�D���HN�G��3�@n��CqCO$8
�;�F��Z3��T0 k� ����2d q51DD"3Q  ��O    �����	�4d�{�D��@N�G�|3�@n��CpCO$8
�7�F��Z3��T0 k� ����2d q51DD"3Q  ��O    �����	�0d�{�D��<N�G�|3�@n��C oCO(7
�7�H���Z3��T0 k� ����2d q51DD"3Q  ��O    �����	�0c�{�D��4N�G�|3�@n��C~�nCO(7
�7�H���Z3��T0 k� ����2d q51DD"3Q ��O    �����	�0c�w�D��,
N�G�|3�@n��C~�mCO,7
�7�H��Z3��T0 k� ����2d q51DD"3Q ��O    �����	�,bw�F�(N�G�|3�E.��C~�mCO,7
�7�H��Z3��T0 k� ����2d q51DD"3Q ��O    �����	�,bw�F�$N�G�|3�E.��C~�lCO06
�7�H��Z3��T0 k� ����2d q51DD"3Q ��O    �����	�,bw�F�$N�G�|3�E.��C~�lCO06
�7�H��Z3��T0 k� ����2d q51DD"3Q ��O    �����	�(aw�F� N�G�|3�E.��CN�kC_46S7�H��Z3��T0 k� ���#�2d q51DD"3Q ��O    �����	�(aw�F� N�G�|3�E.��CN�jC_45S7�H��Z3��T0 k� �#��'�2d q51DD"3Q ��O    ������$`w�F�N�K�|7�E��CN�jC_85S7�H��Z3��T0 k� �'��+�2d q51DD"3Q ��O    ������$_s�F�N�K�|7�E��CN�iC_<5S7�H��Z3��T0 k� �+��/�2d q51DD"3Q  ��O    ������ ^s�F��N�K�|7�E��CN�hC_<4S;�H��Z3��T0 k� �+��/�2d q51DD"3Q  ��O    ������ ^s�F��N�K�|7�E��CN�fC_@4
�;�H��Z3��T0 k� �/��3�2d q51DD"3Q  ��O    ������]o�D���N�K�|;�E��CN�eC_@4
�;�H��Z3��T0 k� �3��7�2d q51DD"3Q  ��O    ������\o�D���N�K�|;�E���CN�cC_D3
�?�H��Z3��T0 k� �7��;�2d q51DD"3Q  ��O    ������\o�D��� N�K�|;�E���CN�bC_D3
�?�H��Z3��T0 k� �7��;�2d q51DD"3Q  ��O    ������[o�D��� N�K�|;�E���CN�`C_H3
�?�H��Z3��T0 k� �;��?�2d q51DD"3Q  ��O    ������Zk�D���� N�K�|;�E���CN�_CoL3
�?�H��Z3��T0 k� �?��C�2d q51DD"3Q  ��O    ������Yg�E~��� N�K�|;�E���E.�]CoL2
�?�H��Z3��T0 k� �<�@2d q51DD"3Q  ��O    ������Xg�E~��� N�K�|;�E���E.�\CoP2
�?�H��Z3��T0 k� �@�D2d q51DD"3Q  ��O    ������V_�E~��� D�K�|?�E�ÒE.�YCoT2
�?�H��Z3��T0 k� �D�H2d q51DD"3Q  ��O    ������U[�E~��� D�O�|?�E�ÒE.�WE�T1
�?�H��Z3��T0 k� �H�L2d q51DD"3Q  ��O    ������S[�E~��� D�O�|?�E�ǒE.�UE�X1
�?�H��Z3��T0 k� �L�P2d q51DD"3Q  ��H    �����oRW�E~��� D�O�|?�E�ǒE.�TE�X0
�?�H��Z3��T0 k� �L�P2d q51DD"3Q  ��H    �����oQ�S�D���� D�O�|?�E�˒E.�RE�\0
�?�H�#�Z3��T0 k� �P�T2d q51DD"3Q  ��H    �����oP�O�D���� D�O�|C�E�˒E.�PE�\/
�?�H�#�Z3��T0 k� �P�T2d q51DD"3Q  ��H    �����oN�K�D���� D�O�|C�E�ϒE.�OE�\/
�?�H�#�Z3��T0 k� �P�T2d q51DD"3Q  ��H    �����oN�C�D�#� l  D�O�|C�E�ӒE.�KE�`.?�H�'�Z3��T0 k� �L�P2d q51DD"3Q  ��H    �����oL�;�F#� l  D�O�|C�E�ӒE.�JE�d-?�H�'�Z3��T0 k� �P�T2d q51DD"3Q  ��H    �����o K�7�F#� l  D�O�|C�E�גE.�HE�d,?�D�+�Z3��T0 k� �P�T2d q51DD"3Q  ��H    �����o I�3�F'� l  D�O�|C�E�ےE.�FAd+;�D�+�Z3��T0 k� �D�H2d q51DD"3Q  ��H    �����n�H�/�F'� l  E�O�|C�E�ےE.�DAd+;�D�+�Z3��T0 k� �<�@2d q51DD"3Q  ��H    �����>�F�'�F+� � E�O�|C�E�ߒE.�CAd*%S;�D�/�Z3��T0 k� �8�<2d q51DD"3Q  ��H    �����>�D�#�F/� � E�O�|@ E��E.�AAd)%S;�D�/�Z3��T0 k� �4�82d q51DD"3Q  ��H    �����>�D��F3� � E�O�|@ E��E.�=Ah'%S7�D�3�Z3��T0 k� �0�42d q51DD"3Q  ��H    �����>�C��D�3� � FS�|@ E��E�;Ad&%S7�D�7�Z3��T0 k� �,�02d q51DD"3Q  ��H    �����>�A��D�7� � FS�|@ B��E�:Ad%%S7�D�7�Z3��T0 k� �,�02d q51DD"3Q  ��H    �����>�?��D�;� � FS�|@ B���E�8Ad%%S7�D�;�Z3��T0 k� �,�02d q51DD"3Q  ��H    �������>���D�;� � FS�|@ B���E�6Ad$%S7�D�?�Z3��T0 k� �(�,2d q51DD"3Q  ��H    �������<���D�?� � FS�|@ B���E�5Ad#%S3�D�?�Z3��T0 k� �(�,2d q51DD"3Q  ��H    �������:���E~?�L D�W�|@ B��E�3Ad"%S3�D�C�Z3��T0 k� �(�,2d q51DD"3Q  ��H    �������:���E~G�L D�W�|@ I�E�0A/`%S3�D�K�Z3��T0 k� �,�02d q51DD"3Q  ��H    �������9���E~G�L 	D�[�|@ I�E�.A/`%S3�D�O�Z3��T0 k� �,�02d q51DD"3Q  ��H    �������7���E~K�L 
D�[�|@ I�E�,A/`%S/�D�O�Z3��T0 k� �,�02d q51DD"3Q  ��H    �������5���E~K�L D�_�|@ I�E�+A/\%S/�D�S�Z3��T0 k� �(	�,	2d q51DD"3Q  ��H    �������3��D�O�L D�_�|@ I�E�)A/\%S/�D�W�Z3��T0 k� �(�,2d q51DD"3Q  ��H    �������1��D�S�L D�c�|@ I/�E��(E?\%S/�D�[�Z3��T0 k� �4�82d q51DD"3Q  ��H    �������/��D�S�L Fc�|@ I/�E��&E?X%S/�D�_�Z3��T0 k� �8�<2d q51DD"3Q  ��H    ������/��D�W�L Fk�|@ I/�E��#E?T%S+�D�g�Z3��T0 k� �<�@2d q51DD"3Q  ��H    ������-��I�W�L Fk�|@ I/�E��"E?T%S+�D�k�Z3��T0 k� �< �@ 2d q51DD"3Q  ��H    ������+��I�[�\Fo�|@ I�E��!E?T%S+�D�o�Z3��T0 k� �C��G�2d q51DD"3Q  ��H    ������)��I�[�\Fs�|@ I�E�� E?P%S+�D�s�Z3��T0 k� �G��K�2d q51DD"3Q  ��H    ������'��I�[�\Fw�|@ I�E��E?P%S+�D�{�Z3��T0 k� �G��K�2d q51DD"3Q  ��H    ������%�I�_�\E�w�|@ I�E��E?P%S+�D��Z3��T0 k� �G��K�2d q51DD"3Q  ��H    ������#w�I�_�\E�{�|@ I#�E��E?L%S'�F��Z3��T0 k� �G��K�2d q51DD"3Q  ��H    ������!o�I�_�,E��|@ I/#�E��E/L%S'�F��Z3��T0 k� �K��O�2d q51DD"3Q  ��H    ������g�I�_�,E���|@ I/#�E~�E/L
%S'�F��Z3��T0 k� �O��S�2d q51DD"3Q  ��H    ����� W�I�_�,!E���|@ I/#�E~�E/H%S'�F��Z3��T0 k� �S��W�2d q51DD"3Q  ��H    ����� K�F_�,"E���|@ I/#�E~�E/H%S'�F��Z3��T0 k� �S��W�2d q51DD"3Q  ��H    ������C�Fc�,$E���|@ I#�E~�E�H%S'�F��Z3��T0 k� �K��O�2d q51DD"3Q  ��H    ������;�Fc�,&E���|@ I#�E~�E�HC'�E���Z3��T0 k� �G��K�2d q51DD"3Q  ��H    ������3�Fc�,(E���|@ I#�E~�E�H C#�E���Z3��T0 k� �C��G�2d q51DD"3Q  ��H    ������+�Fc�,*E���|@ I#�E~�E�G�C#�E���Z3��T0 k� �;��?�2d q51DD"3Q  ��H    ������#�Fg��+E���|@ I#�D��E�G�C#�E���Z3��T0 k� �;��?�2d q51DD"3Q  ��H    �������Fd �-E���|@ @#�D��E�G�C#�E���Z3��T0 k� �;��?�2d q51DD"3Q  ��H    ��������Fd�/E���|@ @#�D��E�G�C#�E���Z3��T0 k� �;��?�2d q51DD"3Q  ��H    ������
��Fh�1E���|@ @#�D��E�G�C#�E���Z3��T0 k� �;��?�2d q51DD"3Q  ��H    ������ ���Fh�3E���|@ @#�D��E�C�C#�E���Z3��T0 k� �7��;�2d q51DD"3Q  ��H    �����                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��� ]�,{,z X �����   + +       ����5    �����l�     b�           ����           � �  �  ���   0		 
 
         ����   � �  ����,    �������       �          V	����         ���     ���    	!
          ��Ȳ          ����    ��Ȳ����                  	����         �     ���  H
          ���s     
    ��1�    ���s��1�                  	����          0     ��� @ 0	 

         ����  � �
	   .��/    �����冉    �� F           R ����           �    ���   @	
          ����  ��	      B�4    �����4                              ���)              �  ���    8

 '            ��B $ $       V�Ȓ�    ��B�Ȓ�                     	    5         ��      ��@   (
 
           kB         j�ۂ�     kB�ۂ�                       v ;         <      ��@   0	
          ���X         ~�{�5    ����{�5    A              	     B          �     ��J   H
D
 
           :�7   �
    � ��     :�� ��     "                �� �         	  �P     ��@   H	$
          l`� � �
      � O��     l] O�[     5                 �         
 [`
`     ��P   03 
          ��O��     � ���    ��O ���                              ���              �  ��@    P		 5                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          +�S  ��        �����     +�L����    �   "                 x                j  �   �   �                          +    ��        ���       +  ��           "                                                �                         ����������������{ � O �������       	 
         
    ��� �J        � �`� � a� �D  ^� �� _  �� 0_@ �  _� �D _� �� d� �� d� �  d����J ����X ����. ����< ����J ����X � � p� �  u� � �r@ �  s@ 
�< V� 
�� V� 
�\ W  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �� �R� � }`���� ����� � �� �j� �� k� �� �o� �� p� �d �[� �d \����� � F� @u@ G u� G$ u� �� `r@ � s  ��  s  � s` B� �m@ 7� `j� 8� @k� � �`� � a� ?� �[� @� 0\� A ]  A$ ]@ 
�\ U� 
�� V  
�| V  
�< V� 
� V� 
� W  
�\ W� 
�� W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������������ e  ������  
�fD
��L���"����D" � j  "  B   J jF�"      �j * , .��
��
��"   "D�j�
�� " �
� �  �  
� ��    ��     ���  �   ����  ��     ���      ��    ��     ��{          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �ODD      ��6 �  ���        � � �  ���        �        ��        �        ��        �    ��    {���p��        ��                         T�) , � ��                                    �                 ����            �������%��  ������                44 Stephane Richer                                                                                  4  3      �`CBi CJ �bCK �k~ � �B� � � B� � �B� � � J� � �	B� � � 
B� � �B� � �B� � � B� � �K � � K � �C � � C" � � �5 � �4 �kV � � k^ � �kjq � kr� �K. � � K6 � � K7 � � K8 � z K9 � r K: � �"� � � "� � � "� � �!*� �""� � #"� �$� � 
� � 
� � � 
� � � 
� � � 
� � �*� � � 
� � ,"P �-!� �=."* |U/"< �] "2 |S !� |P2"< �X "2 | �4� �5
� �  "P � � 7" z �  "E r �  "E r �  "E r � ;" z �  "E rP  *CVP  *CV � )�t                                                                                                                                                                                                                         �� P         �     @ 
        �     i P E j  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    �~�{� ��������������������������������������������������������   �4, d   < s  � �� Ђ�*��0���������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       O    $     �  0$�J      	                             ������������������������������������������������������                                                                                                                                       �    ���                      ��                  
   �� ����� � �������  �� �������������������������� ������� �������������� �  ���� ������������������ �� ��� ������� ��� ��� ��� ���� ���� ���  ���������������������������  ������������������  ������� �������������������� ����������� ���                                     
  5        D��J      �                             ������������������������������������������������������                                                                                                                                        �     s��                      �  �            
 	    ������ � ������������� ����� ���������� �� �� ������������������ ������������������������������ ����� ������  �������� ������� ������� ������������� �������������� ����� ���� ��������������������  �� �������������� �����                                                                                                                                                                                                                                                                                     	                   
                   �             


             �  }�           N                c�                                   �  B                     ����������������  u.  U�    ��������������������������������������������  �����  #&��������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 8 F <                                  � ]7�� �\                                                                                                                                                                                                                                                                                     E)n�  �        m      m                              m      e                                                                                                                                                                                                                                                                                                                                                                                                          
 �  >�  (�  (�  (�  Bm ��
�2 �V ��K����H�+����2��� �����������                ���  � v         �   & AG� �   �                 �                                                                                                                                                                                                                                                                                                                                        7 H   �         #             !��                                                                                                                                                                                                                            Y   �� �� ����      �� v      �� ����� � �������  �� �������������������������� ������� �������������� �  ���� ������������������ �� ��� ������� ��� ��� ��� ���� ���� ���  ���������������������������  ������������������  ������� �������������������� ����������� ��������� � ������������� ����� ���������� �� �� ������������������ ������������������������������ ����� ������  �������� ������� ������� ������������� �������������� ����� ���� ��������������������  �� �������������� �����             "fffffffffffffffffffffffffffffffffffffffffffffff�ff�UflUUfkUUfjWyfffkfffƸww�UUUUuWUuUUUWuUU��UZw��fffl�f��u�UUUYUw�uwwWwUuuWUWWwffffffffffffffff�fffW�ffU�ffUXffffffffffffffffffffffffffffflfffifg��j��ue�uueUUW�Uuw�uUUUuuUWX�U�XuUUXUUUuUUUUUXUW\{U\V�U\{�U[��uwuuUUUWUw���W�XeUl�eUʚeUuU�WWwuU�fWUWf��u���Uv�̅�����UWU�ww��fffff�fffffffff�fffffff�fffffffffffifffhfffhfffiffflffffffffffffYW�UXUWWUUuuUX�U��gUe�kWe��ug���uUUUwWuUUUUUUU��UZf�U\iWUV�xu\��Uww�UUUww���ffff�ffk�fl��ff���f����ux��[����fff��ff��f���f��Vf��fffffffflfff��ff���f̼������˼��jVW�fYY�f���f��wf��xf�yXfiV�fl\kU\wxU�WU��Ww�{ww�{x��|Wx�{wx�{Xxx�hWw��Ww��wx��w����xwzw�x��wx�yWj|�U�Z�uz��u[�yu���x���j�vy���[k���˻��k���l���l���l���l���k̼�ffffffffffffffffffflfff�fff�ff̼ffwilƥ�ffgUl�fuf�Ʃl̶�l��u���W��X�UjXx\hwwyʇw���wuviWy�l�x���w�uXww�x�x��wZ�fw�x�w�x�w���x�x�f��V���ƻ�klf�l�ʉfl�\fl��flh�ff���˼�̻�����̼�������̼�����˼�fl���̼���˻̼�����ƻ�ffffffffff���W��ux��W��uW�eUw��Uw��Ww��Uwxw�ykwy��wu�ywW���u��wwZ���x�w�x���x������ʻ�������̺��ƪ��ƺ��ƻ�ffl�ff̶fflffflfffffff�fffkff̹̻��̻���˻�̻��l˻��˻���˻wx��fffffffffflf�fffffflf��fffffffffffflfffffffffff�ffff�ff�ffffffffI7.    3      A   &�  +                       X     �  �����J���J      ��     �      �   �   �               �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �� ��  � ��     � ��   	 ��   p �� �� ��  � ��  � ��   ��T  ���c@ �� �� �z�c@ AD �$ ��  ��  �� ��   � �� ��     &    { ���8�������J JV<   &    ��  �� �� �  �� �� �z � ��� �$  � �  �� �  �      �  ��   �������2����   g��� 	 �     f ^�         �� !��            ���~���2�������J���j���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                                         �� �����虙������(��������������񙙘�!                �  �������                           �       �  "(� """ �"" ""  "   �      �   �"��"""�"""�"""�"""�����������������������������������""�".�"/��"���!���.���/���-���""����������.���-������/�������   ��  �  .� /�� "�� "� "-�                                ""�  �(��""! ("" �"  �"   ����������������陙����.��� 陙/���.���"���"!��"��".���!♒""����������������̎���""�""",""/ �-� /� "�� "�� . /� �                    �                                           ""陂".��""� � �          �"(��(""������� ��        ""!�"!������������           ��     �                       wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                               s   D   O   w   w   v   u   f   T   �   �              3@  DDp ��4 ��tp��wpO�tpdfwGfeTwfeWwfUFwdUFweTfp�DDp���p���@�w�p   C   D   O   D   w   u   U   U  F  d  f   f   D   �   �   �DD ���7���uP��e`O�V ffg ffG Ufw UU� FUN dFw ffp DDp ��p ��@ w�p  C4 4D@O�C���O�Dt�GVfeVfdFfdFfdUfffUfffwFff�DDD���� ���                    0   G   W   W   U   E   E   w   �   �   @    fg D� O�� �� w�}�w��}����������M���M���M��������y�                    �   �   �   �   �   �   �   �   ~   w       ���w���w���~���~�DMw�������������y�                        w���w}��wt��wt��w}M�����������   M   M   ~�  p�  p   p   p      �   �   �   �               vd  eVp ffpw�Op���w���G���M�}�                                     v   ub  ub  f   `   P               "  f  U` wfP        p   p   p   p   p   p   p   p                               C4 �y�                              f  vU`vf`D�O������p}�w�  ?�  ?�  ?�  33  3#                                      f  Ug	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 " ""   ""     " ""   "" "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "!  "" "  """ !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �            " ""   ""     " ""   "" "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                             �   �   �   �  
� 	�� �� ���	���
���	������+�ݼ� �  
C  �U  �T 
UC 
UT ED  �D  ��  �  �   " �"  �     �        �   ��  ��  ��  w�  ��  ��� ��� ̻� ̻���˩�̽��̽� ˉ� ��  340 UT0 DD0 330 33  C  C  
�  �  ,�  ""  "  �� ��     �      �   ��  �  ��  �             �  �   �   ��  �                                        ��                   �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                                                                                                                                                                
���	���̜̽�˽�̈ۻ��ۻ�۽��˲"������"���" ��"                "   "   "                 ���       �   �  �  ����           �  ��� ݼ� w�� m}� ggp wz�����""H�""T�B"UJ�"UJ�@T�DT�TUJ�  ��.�                           5J� �J� �˻ �˰ ʘ� ̪ ˲"�" ""�"" �  ��                /���"/�  ��                    �                                                                            �               �  �  ��  �   �   �                    �  �˰ ��� �wp ���                                                                                                                                                                �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �   �   �                .                �  �� �� �� ��                         ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                                  �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                                    �   �   �                "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                    �     �                                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                          �  �  �  �� ݚ� }�Ȫ��˙������˼� ��  ��  ��  ��  ��  I� H� �E X�T X�S T�D �[ ˻  ˸  ��  
� �,"��"" "  �" �  ""� �� ˻ �˻ ��ݪ��کɨ��ˀ�̽ ��� ��  ̽  ̻  ̻  ˉ  ��  �D  DC  C3  #;  ;�� �� ��  �� "�  "  �"/ / ����� ��  �      �   �          �  �  "     "  "  "   "�  �  �   �   
                            �          �   �          �                    ��  ���� ��    �����                                             ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                          �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �                    �          �         �   �  �  �   �               �   �               � � ����� ��                                                                                                                                                                                        �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �    �  �   �   ��  �                        �   ������  ��   "   "   "  �� ��                   ����������                                ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                  �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �  "������"    /   �  �   ��                             �                        ���� ��� ����                � ��                    ���� �                             � �������������  �                                 ����                  �   �� �       �  �  ��  �   �   �   �                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �           �  �   �   ��  �                   "   "   "                                   �   �                      �������  ���    �                    ��� ���� ��                   � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        �   ���������  ��            +"  "   " ��������            �� ̽ ̽ ۽�}ک z�� ���๜����̼�ͼ���� �ͼ ��      	            �̀ �ɨ �����ؼ��ݼ ̽� ��� �˰ �˘ ������UP��UZ�UUJ             �                            �   �    �   �     ET DD 
33  33  3       �   DU� UU� ET@ 5[� �ɀ ؚ� ��� +�    �   �                                �   �       �    �                     �   �  �  �    �  �  ��  �   �   �                          � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                           �  �  �  �  �� 
�w ��p������˚��̸���̽��̍̽��̽�����̘�������J�ST�C UJ� Z�  J�  ۼ �� ʨ "�� "+� "" �""   ���   ��  ��  �p  }`  g`  w                   �   �   �   �   �   �   ""  "   ". 0  �@  �   �   �               "�  "/  ����  �       �       �        ���                    ������������                        �                      �                        ���� ��� ����                            ��  ��  ���              �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                                           �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �               � � ����� ��                                                                                                                                                                                               �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""��������D�M����""""�������D�M�M""""�����AMAD������""""��������D��""""������MM�����""""���������D�""""������������������""""������������������������"""$���4���4���4���4���4���4ffffffffffffffffff333DDDffffffffffffffffffffffff3333DDDDafaafffaffDDffff3333DDDDfFfFDfFFfFffdFffff3333DDDDfaffaffaffafffDfffff3333DDDDADAFaFadFfDffff3333DDDDafffDfdFdffff3333DDDDDDFFDfFFfdFffff3333DDDDAffAffaffafffDffffff3333DDDDffffffffffffffffffffffff3333DDDDfff4fff4fff4fff4fff4fff43334DDDD"""������������������""""������������������������""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""���������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��������������D�����3333DDDDI����D��DI����3333DDDDADAIA����D������3333DDDD��������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq`CBi CJ �bCK �k~ � �B� � � B� � �B� � � J� � �	B� � � 
B� � �B� � �B� � � B� � �K � � K � �C � � C" � � �5 � �4 �kV � � k^ � �kjq � kr� �K. � � K6 � � K7 � � K8 � z K9 � r K: � �"� � � "� � � "� � �!*� �""� � #"� �$� � 
� � 
� � � 
� � � 
� � � 
� � �*� � � 
� � ,"P �-!� �=."* |U/"< �] "2 |S !� |P2"< �X "2 | �4� �5
� �  "P � � 7" z �  "E r �  "E r �  "E r � ;" z �  "E rP  *CVP  *CV � )�t3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������.�G�R�K��2�G�]�K�X�I�N�[�Q� � � � � � ��=�@�����������������������������������������!��,�X�K�Z�Z��2�[�R�R� � � � � � � � � � ��=�@�������������������������������������������<�Z�K�V�N�G�T�K��;�O�I�N�K�X� � � � � �=��;�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������=��;� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ������������������=�@� ��!������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            