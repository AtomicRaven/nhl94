GST@�                                                            \     �                                               G  �                        ���������	 J���������������z���        �h      #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"      �j* , . ���
��
�"   "D�j��
� " ��
  d                                                                               ����������������������������������      ��    bbo QQ g 11 44               		� 

                      ��                      nn� ))         888�����������������������������������������������������������������������������������������������������������������������������o=  0  o4   1  +      '           �                    	�  7�  V�  	�                    
          : �����������������������������������������������������������������������������                                �  5     %�   @  #   �   �                                                                                '       )n)n�  
    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�9O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E } �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��o.�_K��P ��2K��q|+� �ץ@�GHm{��\gA��qY�lT0 k� �t�x2d q&�1D"3Q ��?    � ����o.�_K��P ��2K��q|+� �צ@�HHm{��\gA��qY�lT0 k� �t�x2d q&�1D"3Q ��?    � ����p.�_K��P ��2K��q|+� �צ@�HHm��\gA��qY�lT0 k� �x�|2d q&�1D"3Q ��?    � ����p.�^K��P ��3K��q|+� �צ@�HHm��\gA��qY�lT0 k� �|��2d q&�1D"3Q ��?   � ����p.�^K��P ��3K��q|+� �צ@�HHm��\hA��qY�lT0 k� ܀��2d q&�1D"3Q ��?    � ����p.�^K��P ��3K��q|+� �צ@�HHm��\hA��qY�lT0 k� ����2d q&�1D"3Q ��?    � ����q.�^K��P ��3K��q|+� �צ@�HHm���\hA��qY�lT0 k� ����2d q&�1D"3Q ��?    � ����q.�^K��P ��3K��q|+� �צ@�HHm���\hA��qY�lT0 k� ����2d q&�1D"3Q ��?    � ����q.�^K��P ��3K��q|+� �צ@�HA����XhA��qY�lT0 k� ����2d q&�1D"3Q ��?    � ����q.�^K��P ��3K��q|+� �צ@�HA����XhA��qY�lT0 k� ����2d q&�1D"3Q ��?    � ����q.�^L�P ��3K��q|+� �צ@�HA����XhA��qa�lT0 k� ���2d q&�1D"3Q ��?    � ����r.�^L�P ��3K��q|+� �צ@�HA����XhA��pa�lT0 k� ���2d q&�1D"3Q ��?    � ����r.�^L�P ��3K��q|+� �צ@�HA����XhA��pa�lT0 k� ���2d q&�1D"3Q  ��?    � ����r.�^L�P ��3K��q|+� �צ@�HA����XhA��pa�lT0 k� �	��	2d q&�1D"3Q  ��?    � ����r.�^L�P ��3K��q|+� �צ@�HA����XhA��pa�lT0 k� �	��	2d q&�1D"3Q  .�?    � ����r.�^L�P ��4K��q|+� �צ@�HA����XhA��pa�lT0 k� �
��
2d q&�1D"3Q  ��?    � ����s.�^L�P ��4K��q|+� �צ@�HA����XhA��pa�lT0 k� �
��
2d q&�1D"3Q  ��?    � ����s.�^L�P ��4K��q|+� �צ@�HA����XhA��pa�lT0 k� �
��
2d q&�1D"3Q  ��?    � ����s.�^L�P ��4K��q|+� �צ@�HA����XhA��pa�lT0 k� ���2d q&�1D"3Q  ��?    � ����s.�^L�P ��4K��q|+� �צ@�HA����XhA��pa�lT0 k� ���2d q&�1D"3Q  ��?    � ����s.�^L�P ��4K��q|+� �צ@�HA����XhA��pa�lT0 k� ���2d q&�1D"3Q ��?    � ����s.�^L�P ��4K��q|+� �ק@�HA����XhA��pY�lT0 k� ���2d q&�1D"3Q ��?    � ����t.�^L�P ��4K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q ��?    � ���t.�^L�P ��4K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q ��?    � ���t.�^L�P ��4K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q ��?    � ���t.�^L�P ��4K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q ��?    � ���t.�^L�P ��4K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q ��?    � ���t.�^L�P ��4K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q ��?    � ����t.�^L�P ��4K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ����t.�^L�P ��4K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ����t.�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ����s.�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ����s.�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ����s.�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ����s.�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ��~�r.�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ��~�r.�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ��~�q.�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ��~�q.�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ����2d q&�1D"3Q  ��?    � ��~�p�^L�P ��5K��q|+� �ק@�HA����XhA��pY�lT0 k� ��� 2d q&�1D"3Q  ��?    � ��~�p�^L�P ��5B��q|+� �ק@�HA����XhA��pY�lT0 k� � �2d q&�1D"3Q  ��?    � ��~�o�^L�P ��5B��q|+� �ק@�HA����XhA��pY�lT0 k� ��2d q&�1D"3Q  ��?    � ��n�n�^L�P ��5B��q|+� �ק@�HA����XhA��pY�lT0 k� ��2d q&�1D"3Q  ��?    � ��n�m�^L�P ��5B��q|+� �ק@�HA����XhA��pY�lT0 k� ��2d q&�1D"3Q  ��?    � ��n�m�^L�P ��5B��q|+� �ק@�HA����XhA��pY�lT0 k� ��2d q&�1D"3Q  ��?    � ��n�l�^L�P ��5E��q|+� �ק@�HA����ThA��pY�lT0 k� ��2d q&�1D"3Q  ��?    � ��n�k�^L�P ��5E��q|+� �ק@�HA����TiA��pY�lT0 k� ��2d q&�1D"3Q  ��?    � ��n�j�^L�P ��5E��q|+� �ק@�HA����TiA��pY�lT0 k� ��2d q&�1D"3Q  ��?    � ��n�i�^L�P ��5E��q|+� �ר@�HA����TiA��pY�lT0 k� �� 2d q&�1D"3Q  ��?    � ��^�h�^L�P ��6E��q|+� �ר@�HA����TiA��pY�lT0 k� � �$2d q&�1D"3Q  ��?    � ��^�g�^L�P ��6E��q|+� �ר@�HA����TiA��pY�lT0 k� �$�(2d q&�1D"3Q  ��?    � ��^�g�^K��P ��6E��q|+� �ר@�HA����TiA��pY�lT0 k� �(�,2d q&�1D"3Q  ��?    � ��^�f�^K��P ��6E��q|+� �ר@�HA����TiA��pY�lT0 k� �(�,2d q&�1D"3Q  ��?    � ��^�e�^K��P ��6E��q|+� �ר@�HA����TiA��pY�lT0 k� �,�02d q&�1D"3Q  ��?    � ����d�^K��P ��6E��p|+� �ר@�HA����TiA��pY�lT0 k� �0�42d q&�1D"3Q  ��?    � ����c�^K��P ��6B��p|+� �ר@�HA����TiA��pY�lT0 k� �4�82d q&�1D"3Q  ��?    � ����b�^K��P ��6B��p|+� �ר@�HA����TiA��pY�lT0 k� �8�<2d q&�1D"3Q  ��?    � ����b��^K��P ��6B��o|+� �ר@�HA����TiA��pY�lT0 k� �<�@2d q&�1D"3Q  ��?    � ����a��^K��P ��6B��o|+� �ר@�IA����TiA��pY�lT0 k� �<�@2d q&�1D"3Q  ��?    � ����`��^K��P ��6B��o|+� �ר@�IA����TiA��pY�lT0 k� �@�D2d q&�1D"3Q  ��?    � ����_��^A�P ��6B��n|+� �ר@�IA����TiA��pY�lT0 k� �D�H2d q&�1D"3Q  ��?    � ����_��^A�P ��6B��n|+� �ר@�IA����TiA��pY�lT0 k� �H�L2d q&�1D"3Q  ��?    � ����_��^A�P ��6K� m|+� �ר@�IA����TiA��pY�lT0 k� �L�P2d q&�1D"3Q  ��?    � ����_��^A�P ��6K�m|+� �ר@�IA����TiA��pY�lT0 k� �P�T2d q&�1D"3Q  ��?    � ����_��^A�P ��6K�l|+� �ר@�IA����TiA��pY�lT0 k� �P�T2d q&�1D"3Q  ��?    � ����_��^A�Pۤ6K�l|+� �ר@�IA����TiA��pY�lT0 k� �T�X2d q&�1D"3Q  ��?    � ����_��^A�Pۤ6K�l|+� �ר@�IA����TiA��pY�lT0 k� �X�\2d q&�1D"3Q  ��?    � ����_��^A�Pۤ6K�k|+� �ר@�IA����TiA��pY�lT0 k� �\�`2d q&�1D"3Q  ��?    � ����_�^A�Pۤ6K�k|+� �ר@�IA����TiA��pY�lT0 k� �`�d2d q&�1D"3Q  ��?    � ����_�^A�Pۤ6K�j|+� �ר@�IA����TiA��pY�lT0 k� �d�h2d q&�1D"3Q  ��?    � ����_�^A�Pۤ6K�j|+� �ר@�IA����TiA��pY�lT0 k� �d�h2d q&�1D"3Q  ��?    � ����_�^A�Pۤ6K�i|+� �ר@�IA����TiA��pY�lT0 k� �h�l2d q&�1D"3Q  ��?    � ����_�^A�Pۤ6K� i|+� �ר@�IA����TiA��pY�lT0 k� �l�p2d q&�1D"3Q  ��?    � ����_�^A�Pۤ7K�$i|+� �ר@�IA����TiA��pY�lT0 k� �p�t2d q&�1D"3Q  ��?    � ���_�^A�Pۤ7K�(h|+� �ר@�IA����TiA��pY�lT0 k� �t�x2d q&�1D"3Q  ��?    � ���_�^A�Pۤ7K�(h|+� �ר@�IA����TiA��pY�lT0 k� �t�x2d q&�1D"3Q  ��?    � ���_�^A�Pۤ7K�,h|+� �ר@�IA����TiA��pY�lT0 k� �x�|2d q&�1D"3Q  ��?    � ���_�^A�Pۤ7K�0g|+� �ר@�IA����TiA��pY�lT0 k� �|��2d q&�1D"3Q  ��?    � ���_�^A�Pۤ7K�0g|+� �ר@�IA����TiA��pY�lT0 k� �� �� 2d q&�1D"3Q  ��?    � ���_�^A�P�7K�4f|+� �ר@�IA����TiA��pY�lT0 k� �� �� 2d q&�1D"3Q  ��?    � ���_�^A�P�7K�8f|+� �ר@�IA����TiA��pY�lT0 k� �� �� 2d q&�1D"3Q  ��?    � ���_�^A�P�7K�8f|+� �ר@�IA����TiA��pY�lT0 k� ��!��!2d q&�1D"3Q  ��?    � ���_�^A�P�7K�<e|+� �ר@�IA����TiA��pY�lT0 k� ��!��!2d q&�1D"3Q  ��?    � ���_�^A�P�7K�@e|+� �ר@�IA����TiA��pY�lT0 k� ��!��!2d q&�1D"3Q  ��?    � ���_�^A�P�7K�@e|+� �ר@�IA����TiA��pY�lT0 k� ��"��"2d q&�1D"3Q  ��?    � ���_�^A�P�7K�De|+� �ר@�IA����TiA��pY�lT0 k� ��"��"2d q&�1D"3Q  ��?    � ���_�^A�P�7K�Dd|+� �ש@�IA����TiA��pY�lT0 k� ��"��"2d q&�1D"3Q  ��?    � ���_^�^A�P�7K�Hd|+� �ש@�IA����TiA��pY�lT0 k� ��#��#2d q&�1D"3Q  ��?    � ��.�_^�^A�P�7K�Ld|+� �ש@�IA����TiA��pY�lT0 k� ��#��#2d q&�1D"3Q  ��?    � ��.�_^�^A�P�7K�Lc|+� �ש@�IA����TiA��pY�lT0 k� ��#��#2d q&�1D"3Q  ��?    � ��.�^^�^A�P�7K�Pc|+� �ש@�IA����TiA��pY�lT0 k� ��$��$2d q&�1D"3Q  ��?    � ��.�^^�^A�P�7K�Pc|+� �ש@�IA����TiA��pY�lT0 k� ��$��$2d q&�1D"3Q  ��?    � ��.�^�^A�P�7K�Tb|+� �ש@�IA����TiA��pY�lT0 k� ��$��$2d q&�1D"3Q  ��?    � ��.�^�^A�P�7K�Xb|+� �ש@�IA����TiA��pY�lT0 k� ��%��%2d q&�1D"3Q  ��?    � ��.�^�^A�P�7K�Xb|+� �ש@�IA����TiA��pY�lT0 k� ��%��%2d q&�1D"3Q  ��?    � ��.�]�^A�P�7K�\b|+� �ש@�IA����TiA��pY�lT0 k� ��%��%2d q&�1D"3Q  ��?    � ��.�]�^A�P�7K�\a|+� �ש@�IA����TiA��pY�lT0 k� ��%��%2d q&�1D"3Q  ��?    � ��.�]�^A�P�7K�`a|+� �ש@�IA����TiA��pY�lT0 k� ��&��&2d q&�1D"3Q  ��?    � ��.�]�^A�O�7K�`a|+� �ש@�IA����TiA��pY�lT0 k� ��&��&2d q&�1D"3Q  ��?    � ��.�]�^A�O�7K�da|+� �ש@�IA����TiA��pY�lT0 k� ��&��&2d q&�1D"3Q  ��?    � ��.�\�^A�O�7K�d`|+� �ש@�IA����TiA��pY�lT0 k� ��'��'2d q&�1D"3Q  ��?    � ��.�\�^A�O�7K�d`|+� �ש@�IA����TiA��pY�lT0 k� ��'��'2d q&�1D"3Q  ��?    � ��.�\��^A�O�7K�d`|+� �ש@�IA����TiA��pY�lT0 k� ��'��'2d q&�1D"3Q  ��?    � ��.�\��^A�O�7K�d`|+� �ש@�IA����TiA��pY�lT0 k� ��(��(2d q&�1D"3Q  ��?    � ��.�\��^A�O�7K�d`|+� �ש@�IA����TiA��pY�lT0 k� ��(��(2d q&�1D"3Q  ��?    � ��.�\��^A�O�7K�d_|+� �ש@�IA����TiA��pY�lT0 k� ��(��(2d q&�1D"3Q  ��?    � ��.�[��^A�O�8K�d_|+� �ש@�IA����TiA��pY�lT0 k� ��)��)2d q&�1D"3Q  ��?    � ��.�[^�^A�O�8K�d_|+� �ש@�IA����TiA��pY�lT0 k� ��)��)2d q&�1D"3Q  ��?    � ��.�[^�^A�O�8K�d_|+� �ש@�IA����TiA��pY�lT0 k� ��)��)2d q&�1D"3Q  ��?    � ��.�[^�^A�O�8K�d_|+� �ש@�IA����TiA��pY�lT0 k� ��*��*2d q&�1D"3Q  ��?    � ��.�[^�^A�O�8K�d_|+� �ש@�IA����TiA��pY�lT0 k� ��*��*2d q&�1D"3Q  ��?    � ��.�[^�^A�O�8K�d_|+� �ש@�IA����TiA��pY�lT0 k� ��*��*2d q&�1D"3Q  ��?    � ��.�[�^A�O�8K�d_|+� �ש@�IA����TiA��pY�lT0 k� ��+��+2d q&�1D"3Q  ��?    � ��.�Z�^A�O�8K�d_|+� �ש@�IA����TiA��pY�lT0 k� ��+��+2d q&�1D"3Q  ��?    � ��.�Z�^A�O�8K�d_!�+� �ש@�IA����TiA��pY�lT0 k� ��+��+2d q&�1D"3Q  ��?    � ��.�Z�^A�O�8K�d_!�+� �ש@�IA����TiA��pY�lT0 k� ��,��,2d q&�1D"3Q  ��?    � ��.�Z�^A�O�8K�d_!�+� �ש@�IA����TiA��pY�lT0 k� ��,��,2d q&�1D"3Q  ��?    � ��.�Z�^A�O�8K�d_!�+� �ש@�IA����TiA��pY�lT0 k� ��,��,2d q&�1D"3Q  ��?    � ��.�Z�^A�O�8K�d_!�+� �ש@�IA����TiA��pY�lT0 k� ��-� -2d q&�1D"3Q  ��?    � ��.�Z�^A�O�8K�d_!�+� �ש@�IA����TiA��pY�lT0 k� � -�-2d q&�1D"3Q  ��?    � ��.�Y�^A�Oۨ8K�d_!�+� �ש@�IA����TiA��pY�lT0 k� �-�-2d q&�1D"3Q  ��?    � ��.�Y�^A�Oۨ8K�d_!�+� �ש@�IA����TiA��pY�lT0 k� �-�-2d q&�1D"3Q  ��?    � ��.�Y�^A�O۬8K�d_!�+� �ש@�IA����TiA��pY�lT0 k� �.�.2d q&�1D"3Q  ��?    � ��.�Y�^A�O۬8B�d_!�+� �ש@�IA����TiA��pY�lT0 k� �.�.2d q&�1D"3Q  ��?    � ��.�Y�^A�O۬8B�d_!�+� �ש@�IA����TiA��pY�lT0 k� �.�.2d q&�1D"3Q  ��?    � ��.�Y�^A�O۬8B�d_|+� �ש@�IA����TiA��pY�lT0 k� �/�/2d q&�1D"3Q  ��?    � ��.�Y.�^A�O ��8B�d^|+� �ש@�IA����TiA��pY�lT0 k� �/�/2d q&�1D"3Q  ��?    � ��.�Y.�^A�O ��8B�d^|+� �ש@�IA����TiA��pY�lT0 k� �/�/2d q&�1D"3Q  ��?    � ��.�X.�^A�O ��8B�d^|+� �ש@�IA����TiA��pY�lT0 k� �0� 02d q&�1D"3Q  ��?    � ���X.�^A�O ��8B�d]|+� �ש@�IA����TiA��pY�lT0 k� �0� 02d q&�1D"3Q  ��?    � ���X.�^A�O ��8B�d]|+� �ש@�IA����TiA��pY�lT0 k� � 0�$02d q&�1D"3Q  ��?    � ���X.�^A�O ��8B�d]|+� �ש@�IA����TiA��pY�lT0 k� �$1�(12d q&�1D"3Q  ��?    � ���X.�^A�O ��8B�d]|+� �ש@�IA����TiA��pY�lT0 k� �(1�,12d q&�1D"3Q  ��?    � ���X.�^A�O ��8B�d]|+� �ש@�IA����TiA��pY�lT0 k� �(1�,12d q&�1D"3Q  ��?    � ���X.�^A�O ��8B�d]|+� �ש@�IA����TiA��pY�lT0 k� �,1�012d q&�1D"3Q  ��?    � ����X.�^A�O ��8Cd]|+� �ש@�IA����TiA��pY�lT0 k� �02�422d q&�1D"3Q  ��?    � ����X.�^A�O ��8Cd]!�+� �ש@�IA����TiA��pY�lT0 k� �02�422d q&�1D"3Q  ��?    � ����X.�^A�O ��8Cd]!�+� �ש@�IA����TiA��pY�lT0 k� �42�822d q&�1D"3Q  ��?    � ����W.�^A�O ��8Cd]!�+� �ש@�IA����TiA��pY�lT0 k� �83�<32d q&�1D"3Q  ��?    � ����W.�^A�O ��8Cd]!�+� �ש@�IA����TiA��pY�lT0 k� �<3�@32d q&�1D"3Q  ��?    � ����W.�^A�O ��8K�d]!�+� �ש@�IA����TiA��pY�lT0 k� �<3�@32d q&�1D"3Q  ��?    � ����W.�_A�O ��8K�d]!�+� �ש@�IA����TiA��pY�lT0 k� �@4�D42d q&�1D"3Q  ��?    � ����W.�_A�O ��8K�d]!�+� �ש@�IA����TiA��pY�lT0 k� �D4�H42d q&�1D"3Q  ��?    � ����W.�_A�O ��8K�d]!�+� �ש@�IA����TiA��pY�lT0 k� �H4�L42d q&�1D"3Q  ��?    � ����W.�_A�O ��8K�d]!�+� �ש@�IA����TiA��pY�lT0 k� �H4�L42d q&�1D"3Q  ��?    � ����V.�_A�O ��8K�d]!�+� �ש@�IA����TiA��pY�lT0 k� �L5�P52d q&�1D"3Q  ��?    � ����V.�_A�O ��8K�d]!�+� �ש@�IA����TiA��pY�lT0 k� �P5�T52d q&�1D"3Q  ��?    � ����V.�_A�O ��8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �P5�T52d q&�1D"3Q  ��?    � ����V.�_A�O ��8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �T6�X62d q&�1D"3Q  ��?    � ����V.�`A�O ��8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �\8�`82d q&�1D"3Q  ��"    � ����U.�`A�O ��8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �`:�d:2d q&�1D"3Q  ��"    � ����U.�`A�O ��8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �d;�h;2d q&�1D"3Q  ��"    � ����U.�`A�O k�8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �d<�h<2d q&�1D"3Q  ��"    � ����U.�`A�O k�8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �d=�h=2d q&�1D"3Q  ��"    � ����T.�`A�O k�8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �d>�h>2d q&�1D"3Q  ��"    � ����T.�aA�O k�8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �d>�h>2d q&�1D"3Q  ��"    � ����T.�aA�O k�8K�d]|+� �ש@�IA����TiA��pY�lT0 k� �d>�h>2d q&�1D"3Q  ��"    � ����T.�aA�O �8K�`]|+� �ש@�IA����TiA��pY�lT0 k� �d>�h>2d q&�1D"3Q  ��"    � ���T.�aA�O �8K�`]|+� �ש@�IA����TiA��pY�lT0 k� �d>�h>2d q&�1D"3Q  ��"    � ���S.�bA�O �8K�`]|+� �ש@�IA����TiA��pY�lT0 k� �d>�h>2d q&�1D"3Q  ��"    � ���S.�bA�O �8K�`]|+� �ש@�IA����TiA��pY�lT0 k� �d>�h>2d q&�1D"3Q  ��"    � ���S.�bA�O �9K�`]|+� �ש@�IA����TiA��pY�lT0 k� �d>�h>2d q&�1D"3Q  ��"    � ���S.�bA�O��9K�`]|+� �ש@�IA����TiA��pY�lT0 k� �d>�h>2d q&�1D"3Q  ��"    � ��^�S.�cA�O��9K�`]|+� �ש@�IA����TiA��pY�lT0 k� �`>�d>2d q&�1D"3Q  ��"    � ����"h1C���S�E`��|+��C��AEB��c��E�G�_�G�T0 k� �� 2d q&�1D"3Q  ��    ��� ����d1C���S�E`��|+��۸C��@C������@cG�_�?�T0 k� ��2d q&�1D"3Q  ��    ��� ����\1E���W�E`��|+��ӸC��?C������@cG�_�;�T0 k� ��2d q&�1D"3Q  ��    ��� ����P1E���TE`��|+��øC��=C�����@cK�_�/�T0 k� ��2d q&�1D"3Q  ��    ��� ����H0E����TE`��|+�ỸC��<C�{����@cK�_�+�T0 k� ��2d q&�1D"3Q  ��    ��� �ø�D0E����TE`��|+�᳷C��;E�{����E�O�_�'�T0 k� ��� 2d q&�1D"3Q  ��    ��� �Ӵ �</E����TE`��|+�	���C��:E�w����E�O�_��T0 k� ����2d q&�1D"3Q  ��    ��� �Ө"�0/E����T
Ea�|+�	���C��8E�s����E�O�_��T0 k� ����2d q&�1D"3Q  �� 	   ��� �Ӥ"�(.E����TEQ�|+�	���C��7E�o����E�O�_��T0 k� ����2d q&�1D"3Q  �� 	   ��� �Ӡ#� -E����TEQ�|+�	���C��6E�k����AS�_��T0 k� ����2d q&�1D"3Q  � 	   ��� �Ә$�-E����PEQ�|+�	���E��5E�k����AS�[��T0 k� ��
��
2d q&�1D"3Q  �� 	   ��� �ӌ&b,E���	�PEQ�|+�As�E��3E�c�ó�AO�[���T0 k� ����2d q&�1D"3Q  �� 	   ��� ~ӄ'b+E��	�LC��|+�Ao�E��2E�_�÷�AO�[���T0 k� ����2d q&�1D"3Q  �� 	   ��� zӀ'a�*E��	�LC�|+�Ag�EҼ1E�[�÷�E�O�[���T0 k� ����2d q&�1D"3Q  �� 	   ��� v�p)a�)E��	�LC�|+�AW�EҰ0E�S�û�E�K�[���T0 k� ����2d q&�1D"3Q  �� 	   ��� r�h*a�(E��	�LC�|+�AO�EҨ/E�O�û�E�K�[���T0 k� ����2d q&�1D"3Q  �� 	   ��� n�d*a�'E��	�LC�|+�AG�EҤ.E�G�û�E�K�[���T0 k� ����2d q&�1D"3Q  �� 	   ��� j�\+a�&E��	�LC�|+�A?�EҜ-E�C����E�G�[���T0 k� �� �� 2d q&�1D"3Q  �� 	   ��� f�T,a�%D1��	�LC�	|+�A7�EҘ,D2?����E�G�[���T0 k� �x"�|"2d q&�1D"3Q  ��    ��� d�D-a�$D1{�	�L"C�|+�A'�E�+D27����E�C�[���T0 k� �d-�h-2d q&�1D"3Q  ��    ��� b�<-Q�#D1s�	�L#C�|+���E�*D2/����E�?�[�� T0 k� �`1�d12d q&�1D"3Q  ��    ��� `�4.Q�"D1o�	�L$C�|+���E�|)D2+����E�?�[�� T0 k� �X4�\42d q&�1D"3Q  ��    ��� ^�,.Q�!D1g�	�L%C�|+���E�t)D2'����E�;�[�� T0 k� �P6�T62d q&�1D"3Q  ��    ��� \�/Q�D1W�	�L'C�|+����E�d(D2����E�7�[�� T0 k� �@7�D72d q&�1D"3Q  ��    ��� Y3/Q�D1O�	�L(C�|+����E�`'D2����E�3�[��T0 k� �<8�@82d q&�1D"3Q  ��    ��� V3/Q�D1G�	�L)C�|+���E�X'D2����E�3�[��T0 k� �48�882d q&�1D"3Q  ��    ��� S3/Q�D1?�	�L*C�|+���A�P'D2����D�/�[��T0 k� �(7�,72d q&�1D"3Q  ��    ��� P2�0QxD17�	�H+C�|+��߿A�H&D2����D�/�[��T0 k� �6� 62d q&�1D"3Q  ��    ��� M2�0QpDA/�	�H,C�|+����A�@&DA�����D�+�[��T0 k� �4�42d q&�1D"3Q  ��    ��� KR�0Q`DA��H-C�|+����A�0&DA����D�'�[��T0 k� �3�32d q&�1D"3Q  ��    ��� HR�0QXDA��H.D|+�п�ER(&DA����D�'�[��T0 k� � -�-2d q&�1D"3Q  ��    ��� ER�0QPDA��D/D |+�з�ER &DA�÷�D�#�[��T0 k� ��)� )2d q&�1D"3Q  ��    ��� BR�0QHDA��D0D �|+�Я�ER&DAۮ÷�D�#�[��T0 k� ��&��&2d q&�1D"3Q  ��    ��� ?R�0Q@D@���@0D � |+�Ч�ER%DA׮ó�D��[��T0 k� ��"��"2d q&�1D"3Q  ��    ��� <R�0Q8D@���@1D �!|+�П�ER%DAϮó�D��[�|T0 k� �� �� 2d q&�1D"3Q  ��    ��� 9R�1Q(D@���83D �#|+�Ћ�EQ�%DAîï�D��[�tT0 k� ����2d q&�1D"3Q  ��    ��� 6�1A D@���83D �$|+�Ѓ�EQ�%DA��ë�D��[�pT0 k� ����2d q&�1D"3Q  ��    ��� 3�1ADP���44D �%|+��{�EQ�%DQ��ë�D��_�lT0 k� ����2d q&�1D"3Q  ��    ��� 0�1ADP���05D �&|+��s�E��%DQ��ç�D��_�hT0 k� ����2d q&�1D"3Q  ��    ��� -�|1A DP���(6D �(|+��c�E��$DQ��ã�D��_�dT0 k� �� �� 2d q&�1D"3Q  ��    ��� *�t1@�DP���$7D�)|+��[�E��$DQ��ӟ�D��_�`T0 k� ��!��!2d q&�1D"3Q  ��    ��� '�l1@�DP��� 7D�*|+��S�EѼ$EᏱӛ�D��^r`T0 k� ��"��"2d q&�1D"3Q  ��    ��� $�d1@�DP���8D�+|+��K�E�$Eᇱӗ�D��^r\T0 k� ��(��(2d q&�1D"3Q  ��    ��� !�P0@�DP���9D�-|+��7�E�$E�w�ӏ�D��^r\T0 k� ��,��,2d q&�1D"3Q  ��    ��� �H0@�DP���:D�.|+��/�E�$E�o�ӈD��^r\T0 k� �t/�x/2d q&�1D"3Q  ��    ��� �@0@�DP���;D�/|+��'�E�$E�g�ӄD��^r\T0 k� �l2�p22d q&�1D"3Q  ��    ��� 280@�D`��;D�0|+�0�A��%E�_�ӀD��^r\T0 k� �`2�d22d q&�1D"3Q  ��    ��� 2000�D`w���<D�1|+�0�A��%E�W��|D��^�\T0 k� �T2�X22d q&�1D"3Q  ��    ��� 2 /0�D`g���<D�2|+�0�A�p%E�G��t
D���^�`T0 k� �D2�H22d q&�1D"3Q  ��    ��� 2/0�D`c���=C��3|+�?��A�d%E�?��pD���^�`T0 k� �82�<22d q&�1D"3Q  ��    ��� R/0�D`[���=C��4|+����A�\&E�7��hD���^�dT0 k� �03�432d q&�1D"3Q  ��    ��� R.0�E�S���=C��5|+����A�T&E�/��dD���^�dT0 k� �(3�,32d q&�1D"3Q  ��    ��� 
Q�.0�E�K���=C�|6|+����A�L&E�'��`D���^�hT0 k� � 3�$32d q&�1D"3Q  ��    ��� Q�.0pE�;���>C�l7|+����A�<'E���TE���^�pT0 k� �4�42d q&�1D"3Q  ��    ��� Q�.0lE�3�?�>C�h8|+����A�4'E���PE���^�t	T0 k� �4�42d q&�1D"3Q  ��    ��� Q�-0dE�+�?�>C�`9|+����A�,'E���LE���^�x	T0 k� ��4� 42d q&�1D"3Q  ��    �����Q�-0\E�#�?�>C�X:|+���A� (E����DE��^�|	T0 k� ��4��42d q&�1D"3Q  ��    �  ����-0TE��?�=C�P:|+���A�(E����@E��^��	T0 k� ��4��42d q&�1D"3Q  ��    �  ����- LE��?�=C�H;|+���A�)D����8E��^��
T0 k� ��5��52d q&�1D"3Q  ��    � ���, @E��?�=C�8=|+����A� *D����,E��	^��
T0 k� ��6��62d q&�1D"3Q  ��    � ���, <E���?�=C�0=|+����EP�*D����(E��^��
T0 k� ��0��02d q&�1D"3Q  ��    � ��Q�, 4E���?�<C�(>|+����EP�*D���� E��^��
T0 k� ��-��-2d q&�1D"3Q  ��    � ��Q�, 0E���?�<C� ?|+���EP�+E`���F�^��T0 k� ��*��*2d q&�1D"3Q  ��    � ��Q�+ (E���?�;C�@|+��w�EP�+E`���F�^��T0 k� ��(��(2d q&�1D"3Q  ��    � ��Q|+  E���?p:C�A|+��g�EP�,E`���!F�^��T0 k� ��&��&2d q&�1D"3Q  ��    � ��Qt+ E���Oh:C� B|+��_�EP�-E`��3"F�^��T0 k� ��&��&2d q&�1D"3Q  ��    � ��Ql+ E���O`9C��B|+��W�EP�-E`��3 #Er�^��T0 k� ��%��%2d q&�1D"3Q  ��    � ��Qd+ E���OX9C��C|+��S�EP�-E`��2�$Er�^��T0 k� ��%��%2d q&�1D"3Q  ��    � ��Q\*E���OP8C��D|+��K�EP�.E`��2�&Er�^��T0 k� ��%��%2d q&�1D"3Q  ��    � ��QT*D���OH7C��D|+��C�EP�.E`��2�'Er�^��T0 k� ��%��%2d q&�1D"3Q  ��    � ��QH*D���O@7D�E|+��;�E@�.D0��2�)Er�^��T0 k� �x#�|#2d q&�1D"3Q  ��    � ��Q8* !D��O05D�F|+��/�E@�/D0{�2�,Er�^��T0 k� �h!�l!2d q&�1D"3Q  ��    � ��Q0)��"D��O(4D�G|+��'�E@�/D0w�2�-D��^��T0 k� �` �d 2d q&�1D"3Q  ��    � ��Q()��#IߘO 3D�G|+���E@x/D0o�2�.D��^��T0 k� �X �\ 2d q&�1D"3Q  ��    � ��Q )��$IߐO2D�H|+���E@p0D0g�2�0D��^��T0 k� �L�P2d q&�1D"3Q  ��    � ���)��%Iߌ_1D�H|+���E@h0D0_�2�1D�� ^��T0 k� �D�H2d q&�1D"3Q  ��    � ���)��&I߈	_0D�I|+���E@`0D0W�B�2D��!^��T0 k� �<�@2d q&�1D"3Q  ��    � ���)��'I߄
^�/D�I|+���E@X0D0O�B�4D��#^��T0 k� �4�82d q&�1D"3Q  ��    � ����(��*I�x^�.D�K|+����E@D0D0C�B�6D��%^��T0 k� �$�(2d q&�1D"3Q  ��    � ����(��+I�t^�-D|K|+���E@<0D0;�B�7D��&^r�T0 k� ��2d q&�1D"3Q  ��' 	   � ����(��,I�p^�,DtL|+���E@40D@3�B�9D��(^r�T0 k� ��2d q&�1D"3Q  ��' 	   � ����(��-I�l^�+DlL|+���E0,0D@+�B�:D��)^sT0 k� ��2d q&�1D"3Q  ��' 	   � ����(��/I�h^�*DdM|+���E0,0D@#�B�;D��*^sT0 k� ��2d q&�1D"3Q  �' 	   � ����(�1E�`^�(DPN|+��תE0$0D@�B�=Er�-^sT0 k� ����2d q&�1D"3Q ��/ 	   � ���'�2E�\n�'DHN|+��ϨE0 0E`�B�>Er�.^s$T0 k� ����2d q&�1D"3Q ��/ 	   � ���'�3E�Xn�%E_@O|+��˦G 0E`�R�?Er�/^s,T0 k� ����2d q&�1D"3Q ��/ 	   � ���'�4E�Tn�$E_8O|+��ǥG 0Eo��R�@Er�1^s4T0 k� ����2d q&�1D"3Q ��/ 	   � ���'�5E�Pn�#E_0P|+����G 1Eo��R�AEr�2^s<T0 k� ����2d q&�1D"3Q ��/ 	   � ���'�6E�Ln�"E_(P|+����G 1Eo��R�BEr�4^sDT0 k� ����2d q&�1D"3Q ��/ 	   � ����'�7E�H�!E_ Q|+����G 1Eo��R�CEr�5^sHT0 k� ����2d q&�1D"3Q ��/ 	   � ��Є'�8FD� E_Q|+����G1Eo��R�DEr�7^�HT0 k� ������2d q&�1D"3Q ��/ 	   � ���t&��:F@�pE_R|+����G1Eo��R�EEr�:^�HT0 k� ������2d q&�1D"3Q ��/ 	   � ���l&��;F<!�hE_ R|+����G 1E_�R�FEr�;^�HT0 k� ������2d q&�1D"3Q ��/ 	   � ���d&��<F8"�`E^�S|+����G�1E_�R�FEb�=^�HT0 k� ������2d q&�1D"3Q ��/ 	   � ���\&��=F4$�XE^�S|+����G/�1E_��|GEb�?YsHT0 k� ������2d q&�1D"3Q �/ 
   � ��PP&��=F4%nPI��T|+����G/�2E_��tGEb�@YsHT0 k� ������2d q&�1D"3Q	 �/ 
   � ��PH&��>F0'nHI��T|+����G/�2E_��pHEb�BYsHT0 k� �����2d q&�1D"3Q	 ��/ 
   � ��P@&��?F0(n@I��T|+����G/�2E_�	�lHEb�DYsHT0 k� �w��{�2d q&�1D"3Q	 ��/ 
   � ��P8&�?F,*n8I��U|+��{�G/�2E_�
�hIEb�EYsHT0 k� �o��s�2d q&�1D"3Q
 ��/ 
   � ��P0%�@F,,n0I��U|+��w�G/�2E_��dIEb�G^�HT0 k� �g��k�2d q&�1D"3Q
 ��/ 
   � ��P(%�@F,-n(I��U|+��o�G/�2E_��`JEb�I^�LT0 k� �[��_�2d q&�1D"3Q
 ��/ 
   � ��@ %�AE�(/n I��U|+��k�G/�2E_��\JEb�J^�LT0 k� �S��W�2d q&�1D"3Q
 ��/ 
   � ��@%�AE�(0^I��U|+��g�G/�2E_|�XKA��L^�LT0 k� �K��O�2d q&�1D"3Q ��/
   � ��@%_�AE�(2^I��U|+��_�G/�2E_t�PKA��M^�LT0 k� �C��G�2d q&�1D"3Q ��/ 
   � ��@%_�BE�(3^I��U|+��[�G/�3E_l�LLA��NY�LT0 k� �;��?�2d q&�1D"3Q ��/ 
   � ��@%_�BE�(5^ I��U|+��W�G/�3E_d�HLA��PY�LT0 k� �3��7�2d q&�1D"3Q ��/ 
   � ����%_�CE�(6]�I��U|+��O�G/�4EO\�DLA��QY�LT0 k� �'��+�2d q&�1D"3Q ��/ 
   � ����%_�CE�(8]�I��U|+��K�G/�4EOT�@MA��SY�LT0 k� ���#�2d q&�1D"3Q ��/    � ����%_�DE�(9]�I��U|+��C�G/�4EOL�@MA��TY�PT0 k� ����2d q&�1D"3Q ��/    � ����%_�DE�(;]�
I��U|+��?�G/�5EOD�<NA��UY�PT0 k� ����2d q&�1D"3Q ��/    � ����%_�EE�(<]�I��U|+��;�G/�5EO<�8NA��WY�PT0 k� ����2d q&�1D"3Q ��/    � ����%_�EE�(=]�I��U|+��3�G/�5C�0�4NA��XY�PT0 k� ������2d q&�1D"3Q ��/   � ����%_�FE�,?]�I��U|+��/�G/�6C�(�0OA��YY�PT0 k� �����2d q&�1D"3Q ��/    � ����%_�FE�,@M�I��U|+��+�G/�6C� �,OA��[Y�PT0 k� ����2d q&�1D"3Q ��/    � ����%o�GE�,AM�I�|U|+��#�@��6C��(PA��\Y�PT0 k� ����2d q&�1D"3Q ��/    � ����%o�GE�0BM�I�xU|+���@��6C��$PA��]Y�PT0 k� �۲�߲2d q&�1D"3Q ��/   � ����&o�HE�0CM�I�tU|+���@��7C�� PA��^Y�PT0 k� �Ӱ�װ2d q&�1D"3Q ��/    � ����&o�HE�0DM�I�tU|+���@��7C���QA��`Y�PT0 k� �ǭ�˭2d q&�1D"3Q
 ��/    � ����&o�HE�4EM�I�pU|+���@��7C���QA��aY�TT0 k� ����ê2d q&�1D"3Q
 ��/    � ����'o�IE�4FM�I�lU|+���@��7C���QA��bY�TT0 k� ������2d q&�1D"3Q
 ��/    � ����'o�IE�8GM�I�lU|+���@��8C�� �RA��cY�TT0 k� ������2d q&�1D"3Q
 ��/    � ����(o�JE�8GMx LhU|+����@��8C�� �RA��dY�TT0 k� ������2d q&�1D"3Q	 ��/    � ���|(o�JE�<HMp LhU|+����@��8C�� �SA��eY�TT0 k� ������2d q&�1D"3Q	 ��/    � ���t)o�KE�<I=g�LdU|+���@��8C��!�SA��fY�TT0 k� ������2d q&�1D"3Q	 ��/    � ���l)o�KE�@I=_�LdU|+���@��9C��!�SA��gY�TT0 k� ������2d q&�1D"3Q ��/    � ���d*o�KE�@J=W�L`U|+���@��9C��!�SA��hY�TT0 k� ������2d q&�1D"3Q ��/    � ���\*o�LE�DJ=O�L`U|+���@��9C��!�TA��iY�T
T0 k� �{���2d q&�1D"3Q ��/    � ���T+o�LE�DK=G�L\U|+��ߎ@��9C��!� TA��jY�T
T0 k� �s��w�2d q&�1D"3Q ��?    � ���L+o�ME�DK�?�L\U|+��ێ@��:EN�!��TA��kY�T
T0 k� �g��k�2d q&�1D"3Q ��?    � ���D,o�ME�HK�7�LXU|+��ӏ@��:EN�!��UA��lY�X
T0 k� �_��c�2d q&�1D"3Q ��?    � ���8-o�ME�HK�/�LXU|+��Ϗ@��:EN�!��UA��mY�X
T0 k� �W��[�2d q&�1D"3Q ��?    � ���0-o�NE�HL�'�LTU|+��ˏ@��:EN�!��UA��nY�X
T0 k� �O��S�2d q&�1D"3Q ��?    � ���(.o�NAHL��LTU|+��Ð@��:ENt!��VA��oY�X
T0 k� �G��K�2d q&�1D"3Q ��?    � ��� /o�NAHL	} LPU|+����@��;ENl!��VA��pY�X
T0 k� �?}�C}2d q&�1D"3Q )�?    � ���/o�OALL	} LPU|+����@��;ENd!��VA��qY�X
T0 k� �3~�7~2d q&�1D"3Q ��?    � ���0o�OALL	} L.LU|+����@��;ENX!��VA��rY�X
T0 k� �+�/2d q&�1D"3Q ��?    � ���1o�OALL	}  L.LU|+����@��;ENP ��WA��sY�X
T0 k� �#�'2d q&�1D"3Q ��?    � ��� 1o�PA_HM	|� L.HU|+����@��;E>H ��WA��tY�X
T0 k� ����2d q&�1D"3Q ��?    � ����2o�PA_HML� L.HU|+����@��<E>< ��WA��uY�X
T0 k� ����2d q&�1D"3Q ��?    � ����3o�PA_HML� L.HU|+����@��<E>4��XA��uY�X
T0 k� ����2d q&�1D"3Q ��?    � ����4o�QA_HML�L.DU|+����@��<E>,��XA��vY�X	T0 k� ����2d q&�1D"3Q ��?    � ����5o�QA_HML�L.DU|+����@�|<E>$��XA��wY�X	T0 k� ������2d q&�1D"3Q ��?    � ����5o�QC�DML�L.@U|+����@�|<E>��XA��xY�\	T0 k� ����2d q&�1D"3Q ��?    � ����6o�RC�DML�L.@U|+����@�x=E>��YA��yY�\	T0 k� ����2d q&�1D"3Q ��?    � ��N�7o�RC�@NL�L.@U|+����@�x=E>��YA��zY�\	T0 k� �߅��2d q&�1D"3Q ��?    � ��N�8o�RC�@NL�L.<U|+����@�t=E> ��YA��zY�\	T0 k� �׆�ۆ2d q&�1D"3Q ��?    � ��N�9o�SC�<NL�L.<U|+���@�t=E=���YA��{Y�\	T0 k� �χ�Ӈ2d q&�1D"3Q  ��?    � ��N�:o�SC�<NL�L.8U|+��w�@�p=E=���YA��|Y�\	T0 k� �ǈ�ˈ2d q&�1D"3Q  ��?    � ��N�;o�SC�8NL�L.8U|+��s�@�p=E-���ZA��}Y�\	T0 k� ��È2d q&�1D"3Q  .�?    � ��N�;o�SC�4NL�L.8U|+��o�@�p>E-���ZA��}Y�\	T0 k� ����2d q&�1D"3Q  ��?    � ��N�<o�TC�4N<�L.4U|+��g�@�l>E-���ZA��~Y�\	T0 k� ������2d q&�1D"3Q  ��?    � ��N�=o�TM0N<�L.4U|+��c�@�l>E-���ZA��Y�\	T0 k� ������2d q&�1D"3Q  ��?    � ��N�>o�TM,O<�L.4U|+��_�@�h>E-���[A��~Y�\	T0 k� ������2d q&�1D"3Q  ��?    � ��>�?o�UM,O<�L.0U|+��[�@�h>E-���[A��~Y�\	T0 k� ������2d q&�1D"3Q  ��?    � ��>|@o�UM(O<�L.0U|+��S�@�h>E-���[A��~Y�\	T0 k� ������2d q&�1D"3Q  ��?    � ��>tA_�UM$O<�L.0U|+��O�@�d>E-���[A��~Y�\	T0 k� �����2d q&�1D"3Q  ��?    � ��>lB_�UM$O<�L.,U|+��K�@�d?E-���[A��}Y�\	T0 k� {���2d q&�1D"3Q  ��?    � ��>dD_�VM O<xL.,U|+��G�@�`?E-���\A��}Y�\	T0 k� s��w�2d q&�1D"3Q  ��?    � ��>\E_�VMO<tL.,U|+��C�@�`?E���\A��}Y�\T0 k� k��o�2d q&�1D"3Q  ��?    � ��>XF_�VMO<l	L.(U|+��;�@�`?E���\A��}Y�`T0 k� c��g�2d q&�1D"3Q  ��?    � ��>PG_�VMP<h
L.(U|+��7�@�\?E���\A��}Y�`T0 k� �[��_�2d q&�1D"3Q  ��?    � ��>PG��VM/P<d
L.$V|+��3�@�\?E���\A��|Y�`T0 k� �S��W�2d q&�1D"3Q  ��?    � ��>LG��WM/P<\L.$V|+��/�@�\?E�
��]A��|Y�`T0 k� �G��K�2d q&�1D"3Q  ��?   � ��>HH��WM/P �XL. W|+��'�@�X@E�	��]A��|Y�`T0 k� �?��C�2d q&�1D"3Q  ��?    � ��.HH��WM/P �TL.X|+��#�@�X@E���]A��|Y�`T0 k� �7��;�2d q&�1D"3Q  ��?    � ��.DI��WM/P �LL.X|+���@�X@E���]A��{Y�`T0 k� �/��3�2d q&�1D"3Q  ��?    � ��.@I��WM/P �HL.Y|+���@�T@E���]A��{Y�`T0 k� �'��+�2d q&�1D"3Q  ��?    � ��.<J��WM/P �DL.Y|+��@�T@@���]A��{Y�`T0 k� ���#�2d q&�1D"3Q  ��?    � ��.<K��WM/P �@L.Z|+��@�T@@���^A��{Y�`T0 k� ����2d q&�1D"3Q  ��?    � ��.8K��WM/P �8L.Z|+��@�P@@���^A��{Y�`T0 k� ����2d q&�1D"3Q  ��?    � ���4L��WM Q �4L.[|+��@�P@@���^A��zY�`T0 k� ����2d q&�1D"3Q  ��?    � ���4M�WM Q �0L.\|+��@�PA@|��^A��zY�`T0 k� �����2d q&�1D"3Q  ��?    � ���0N�WM�Q �,L.\|+���@�LA@x ��^A��zY�`T0 k� ������2d q&�1D"3Q  ��?    � ���0N�WM�Q �(L.]|+���@�LA@w���^A��zY�`T0 k� ����2d q&�1D"3Q  $�?    � ���,O�WM�Q �$L.]|+���@�LA@s���_A��zY�`T0 k� ����2d q&�1D"3Q  ��?    � ���,P�WM�Q �L.^|+����@�LA@o���_A��zY�`T0 k� ����2d q&�1D"3Q  ��?    � ���(P�WM�Q �L ^|+���@�HA@o���_A��yY�`T0 k� ����2d q&�1D"3Q  ��?    � ���(P�WM�Q �L�_|+���@�HA@k���_A��yY�`T0 k� ����2d q&�1D"3Q  ��?    � ���(P�WM�Q �L�_|+���@�HA@g���_A��yY�`T0 k� ����2d q&�1D"3Q  ��?    � ���$Q�WC��Q �L�`|+���@�HA@c���_A��yY�`T0 k� ����2d q&�1D"3Q  ��?    � ���$Q�WC��Q �L�`|+���@�DB@_���_A��yY�dT0 k� ����2d q&�1D"3Q  ��?    � ���$R�WC��Q �L�a|+���@�DB@_���`A��yY�dT0 k� ����2d q&�1D"3Q  ��?    � ��� S�XC��R � L�a|+���@�DB@[���`A��xY�dT0 k� ����2d q&�1D"3Q  ��?    � ��� S��XC��R ��L�a|+���@�@B@W���`A��xY�dT0 k� ����2d q&�1D"3Q  ��?    � ���T��XC��R ��L�b|+���@�@B@W���`A��xY�dT0 k� ����2d q&�1D"3Q  ��?    � ���T��XC��R ��L�b|+���@�@B@S���`A��xY�dT0 k� ����2d q&�1D"3Q  ��?    � ���U��XC��R ��L�b|+� l�@�@B@O���`A��xY�dT0 k� ����2d q&�1D"3Q  ��6    � ���U��XC��R ��L�c|+� l�@�@B@K���`A��xY�dT0 k� ����2d q&�1D"3Q  ��6    � ���V�|XC��R ��L�c|+� lߘ@�<B@K���`A��xY�dT0 k� �����2d q&�1D"3Q  ��6    � ���V�xXC��R ��L�c|+� lߘ@�<B@G���aA��wY�dT0 k� �����2d q&�1D"3Q  ��6    � ���W�tXC��R ��L�d|+� lߘ@�<B@C���aA��wY�dT0 k� �����2d q&�1D"3Q  ��6    � ���W�pXC��R ��L�d|+� �ߘ@�<C@C���aA��wY�dT0 k� ����2d q&�1D"3Q  ��6    � ���W�lXC��R ��L�d|+� �ߘ@�8C@?���aA��wY�dT0 k� ����2d q&�1D"3Q  ��6    � ���W�hXC��R ��L�e|+� �ߘ@�8C@?���aA��wY�dT0 k� ����2d q&�1D"3Q  �6    � ���WdXC��R ��L�e|+� �ߙ@�8C@;���aA��wY�dT0 k� ������2d q&�1D"3Q  ��?    � ���X`XC��R ��L�e!�+� �ߙ@�8C@7���aA��wY�dT0 k� �����2d q&�1D"3Q  ��?    � ���XXXC��R ��L�f!�+�ߙ@�8C@7���aA��vY�dT0 k� ����2d q&�1D"3Q  ��?    � ���XTXC��R ��L�f!�+�ߙ@�4C@3���bA��vY�dT0 k� ����2d q&�1D"3Q  ��?    � ���YPXC��R ��L�f!�+�ߚ@�4C@3���bA��vY�dT0 k� ���#�2d q&�1D"3Q  ��?    � ���YHXC��R ��L�f!�+�ߚ@�4C@/���bA��vY�dT0 k� �'��+�2d q&�1D"3Q  ��?    � ���YDXC��R ��L-�g!�+�ߚ@�4C@/���bA��vY�dT0 k� �/��3�2d q&�1D"3Q  ��?    � ���Z@XC��R ��L-�g!�+��ߚ@�4C@+���bA��vY�dT0 k� �;��?�2d q&�1D"3Q  ��?    � ���Z8XD�R �� L-�g!�+��ߛ@�0C@'���bA��vY�dT0 k� �C��G�2d q&�1D"3Q  ��?    � ��� Z4XD�R �� L-�h!�+��ߛ@�0D@'���bA��vY�dT0 k� �O��S�2d q&�1D"3Q  ��?    � ��� [,XD�R �� L-�h!�+��ߛ@�0D@#���bA��vY�dT0 k� �W��[�2d q&�1D"3Q  ��?   � ��� [$XD�R ��!L-�h!�+��ߛ@�0D@#���bA��uY�dT0 k� �c��g�2d q&�1D"3Q  �?    � ��� [ XD�R ��!L-�h|+��ߛ@�0D@���bA��uY�dT0 k� -_��c�2d q&�1D"3Q  ��?    � ����\XD�R ��"L-�i|+��ߜ@�0D@���cA��uY�dT0 k� -[��_�2d q&�1D"3Q  ��?    � ����\YD�R ��"L-�i|+��ߜ@�,D@���cA��uY�hT0 k� -W��[�2d q&�1D"3Q  ��?    � ����\YD�R۬"L-�i|+��ߜ@�,D@��|cA��uY�hT0 k� -S��W�2d q&�1D"3Q  ��?    � ����]YD�Rۨ#L-�j|+��ۜ@�,D@��|cA��uY�hT0 k� -O��S�2d q&�1D"3Q  ��?    � ����]�YD�Rۨ#L-�j|+��ۜ@�,D@��|cA��uY�hT0 k� �O��S�2d q&�1D"3Q  ��?    � ����]�YD�Rۤ#L-�j|+��۝@�,D@��|cA��uY�hT0 k� �K��O�2d q&�1D"3Q  ��?    � ����]�YD�Rۤ#L-�j|+��۝@�,D@��|cA��uY�hT0 k� �G��K�2d q&�1D"3Q  ��?    � ����^�YD�R۠$L-�k|+��۝@�,D@��|cA��uY�hT0 k� �K��O�2d q&�1D"3Q  ��8    � ����^�YD�Rۜ$L-�k|+��۝@�(DE���xcA��tY�hT0 k� �C��G�2d q&�1D"3Q  ��8    � ����^	��YD�Rۜ$L-�k|+��۝@�(DE���xcA��tY�hT0 k� �7��;�2d q&�1D"3Q  ��8    � ����^	��YD�Rۘ%L-�k!�+��۝@�(DE���xcA��tY�hT0 k� �3��7�2d q&�1D"3Q  ��8    � ����_	��YA�Qۘ%L-�l!�+��۞@�(EE���xcA��tY�hT0 k� �/��3�2d q&�1D"3Q  ��8    � ����_	��ZA�Q۔%L-�l!�+��۞@�(EE���xdA��tY�hT0 k� �+��/�2d q&�1D"3Q  ��8    � ����_	��ZA�Q۔&L-�l!�+��۞@�(EE���xdA��tY�hT0 k� �+��/�2d q&�1D"3Q  ��8    � ����_	��ZA�Qې&L-�l!�+��۞@�(EE���tdA��tY�hT0 k� �+��/�2d q&�1D"3Q  ��8    � ����`	��ZA�Qې&L-�l!�+��۞@�$EE���tdA��tY�hT0 k� �+��/�2d q&�1D"3Q  ��8    � ����`	��ZA�Q�&L-�m!�+��۞@�$EE���tdA��tY�hT0 k� �+��/�2d q&�1D"3Q  ��8    � ����`	��[A�Q�'L-�m!�+��۟@�$EE���tdA��tY�hT0 k� �+��/�2d q&�1D"3Q  ��8    � ����`	��[A�Q�'L-�m!�+��۟@�$EE��tdA��tY�hT0 k� �'��+�2d q&�1D"3Q  ��8    � ����a	��[A�Q�'L-�m!�+� �۟@�$EE��tdA��tY�hT0 k� �#��'�2d q&�1D"3Q  ��8    � ����a	��[A�Q�'L-�m!�+� �۟@�$EE��tdA��tY�hT0 k� �#��'�2d q&�1D"3Q  ��8    � ����a	��[A�Q�(L-�n|+� �۟@�$EE��pdA��sY�hT0 k� �#��'�2d q&�1D"3Q  ��8    � ����a	��[A�Q�(L-�n|+� �۟@�$EE��pdA��sY�hT0 k� �#��'�2d q&�1D"3Q  ��8    � ����b	��[A�Q�(L-�n|+� �۟@� EE���pdA��sY�hT0 k� �#��'�2d q&�1D"3Q  ��8    � �� m�b	��[A�Q�|(L-�n|+� �۠@� EE���pdA��sY�hT0 k� �'��+�2d q&�1D"3Q  ��8    � �� m�b��[A�Q�|)L-�n|+� �۠@� EE���peA��sY�hT0 k� �'��+�2d q&�1D"3Q  ��8    � �� m�b��[A�Q�|)L-�o|+� �۠@� EE���peA��sY�hT0 k� �+��/�2d q&�1D"3Q  ��8    � �� m�c��[A�Q�x)L-�o|+� �۠@� EE���peA��sY�hT0 k� �+��/�2d q&�1D"3Q  ��8    � �� m�c��[A�Q�x)L-�o|+� �۠@� EE���leA��sY�hT0 k� �/��3�2d q&�1D"3Q  ��8    � ����c��\A�Q�t*L-�o|+� �۠@� EE}��leA��sY�hT0 k� �/��3�2d q&�1D"3Q  ��8    � ����c�\A�Q�t*L-�o|+� �۠@� FE}#��leA��sY�hT0 k� �/��3�2d q&�1D"3Q  ��8    � ����c�\A�Q�t*L-�o|+� �ۡ@� FE}#��leA��sY�hT0 k� �3��7�2d q&�1D"3Q  ��8    � ����d�\A�P�p*L-�p|+� �ۡ@�FE}'��leA��sY�hT0 k� �3��7�2d q&�1D"3Q  ��8    � ����d��]A�P�l+L-�p|+� �ۡ@�FH�+��leA��sY�hT0 k� �/��3�2d q&�1D"3Q  ��8    � ����d��]A�P�l+L�p|+� �ۡ@�FH�/��leA��sY�hT0 k� �'��+�2d q&�1D"3Q  ��8    � ����e��]A�P�l+L�p|+� �ۡ@�FH�/��leA��sY�hT0 k� �#��'�2d q&�1D"3Q  ��8    � ����e��^A�P�h+L�p|+� �ۡ@�FH�3��heA��rY�hT0 k� ���#�2d q&�1D"3Q  ��8    � ����e��^A�P�l+L�q|+� �ۡ@�FH�3��heA��rY�hT0 k� ���#�2d q&�1D"3Q  ��8    � ����e��^A�P�l,L�q|+� �ۡ@�FH�7��heA��rY�hT0 k� ����2d q&�1D"3Q  ��8    � ��� e��^A�P�l,L�q|+� �ۢ@�FH�7��heA��rY�hT0 k� ����2d q&�1D"3Q  ��8    � ���f��^A�P�l,L�q|+� �ۢ@�FH�;��heA��rY�lT0 k� ����2d q&�1D"3Q  ��8    � ���f��^A�P�p,L�q|+� �ۢ@�FH�;��hfA��rY�lT0 k� ���#�2d q&�1D"3Q  ��8    � ���f��^A�P�p,L�q|+� �ۢ@�FH�?��hfA��rY�lT0 k� ���#�2d q&�1D"3Q  ��8   � ���f�^A�P�p-L�q|+� �ۢ@�FH�?��hfA��rY�lT0 k� �#��'�2d q&�1D"3Q  ��8    � ��f�^A�P�p-A]�q|+� �ע@�FH�C��hfA��rY�lT0 k� �#��'�2d q&�1D"3Q  ��8    � ��g�^A�P�p-A]�q|+� �ע@�FH�C��hfA��rY�lT0 k� �'��+�2d q&�1D"3Q  ��8    � ��g�^A�P�t-A]�q|+� �ע@�FH�C��dfA��rY�lT0 k� �'��+�2d q&�1D"3Q  ��8    � �� g�^A�P�t-A]�q|+� �ע@�FH�G��dfA��rY�lT0 k� �+��/�2d q&�1D"3Q  ��8   � ��$g�^A�P�t-A]�q|+� �ף@�FH�G��dfA��rY�lT0 k� �+��/�2d q&�1D"3Q  ��8    � ���,g�^A�P�t.A��q|+� �ף@�FH�K��dfA��rY�lT0 k� �+��/�2d q&�1D"3Q  ��8    � ���0g�^A�P�x.A��q|+� �ף@�FH�K��dfA��rY�lT0 k� �/��3�2d q&�1D"3Q  ��8    � ���4h�^A�P�x.A��q|+� �ף@�FH�O��dfA��rY�lT0 k� �/��3�2d q&�1D"3Q  ��8    � ���8h�^A�P�x.A��q|+� �ף@�FH�O��dfA��rY�lT0 k� �3��7�2d q&�1D"3Q  ��8    � ���<h�^A�P�x.A��q|+� �ף@�FH�O��dfA��rY�lT0 k� �3��7�2d q&�1D"3Q  ��8    � ���@h�^A�P�x.A��q|+� �ף@�GH�S��dfA��rY�lT0 k� �7��;�2d q&�1D"3Q  ��8    � ���Dh�^A�P�|.A��q|+� �ף@�GH�S��dfA��rY�lT0 k� �7��;�2d q&�1D"3Q  ��8    � ���Hh�^A�P�|/A��q|+� �ף@�GH�W��dfA��rY�lT0 k� �7��;�2d q&�1D"3Q  ��8    � ���Li�_A�P�|/A��q|+� �ף@�GH�W��dfA��rY�lT0 k� �;��?�2d q&�1D"3Q  ��8    � ���Ti�_A�P�|/A��q|+� �ף@�GH�W��`fA��qY�lT0 k� �;��?�2d q&�1D"3Q  ��8    � ���Xi�_A�P�|/BM�q|+� �פ@�GH�[��`fA��qY�lT0 k� �;��?�2d q&�1D"3Q  ��8    � ���\i�_A�P�|/BM�q|+� �פ@�GH�[��`fA��qY�lT0 k� �?��C�2d q&�1D"3Q  ��8    � ���`i�_A�Pۀ/BM�q|+� �פ@�GH�[��`fA��qY�lT0 k� �?��C�2d q&�1D"3Q  ��8    � ���di�_A�P ��/BM�q|+� �פ@�GH�_��`gA��qY�lT0 k� �C��G�2d q&�1D"3Q  ��8    � ���di�_A�P ��0BM�q|+� �פ@�GH�_��`gA��qY�lT0 k� �C��G�2d q&�1D"3Q  ��8    � ���hj�_A�P ��0B��q|+� �פ@�GH�c��`gA��qY�lT0 k� �C��G�2d q&�1D"3Q  ��8    � ���lj�_A�P ��0B��q|+� �פ@�GH�c��`gA��qY�lT0 k� �G��K�2d q&�1D"3Q  ��8    � ���pj�_A�P ��0B��q|+� �פ@�GH�c��`gA��qY�lT0 k� �G��K�2d q&�1D"3Q  ��8    � ���tj�_A�P ��0B��q|+� �פ@�GH�g��`gA��qY�lT0 k� �G��K�2d q&�1D"3Q  ��8   � ���tj�_A�P ��0B��q|+� �פ@�GH�g��`gA��qY�lT0 k� �7��;�2d q&�1D"3Q  �8    � ���tj�_A�P ��0K��q|+� �פ@�GH}g��`gA��qY�lT0 k� �'��+�2d q&�1D"3Q ��?    � ���tk�_A�P ��0K��q|+� �פ@�GH}g��`gA��qY�lT0 k� ����2d q&�1D"3Q ��?    � ���xk�_A�P ��1K��q|+� �פ@�GH}k��`gA��qY�lT0 k� ����2d q&�1D"3Q ��?    � ���xk�_A�P ��1K��q|+� �ץ@�GH}k��`gA��qY�lT0 k� ������2d q&�1D"3Q ��?    � ���|l�_A�P ��1K��q|+� �ץ@�GH}k��`gA��qY�lT0 k� ������2d q&�1D"3Q ��?    � ���|l�_A�P ��1K��q|+� �ץ@�GHmo��\gA��qY�lT0 k� ������2d q&�1D"3Q ��?   � ����l�_A�P ��1K��q|+� �ץ@�GHmo��\gA��qa�lT0 k� ������2d q&�1D"3Q ��?    � ����l�_A�P ��1K��q|+� �ץ@�GHmo��\gA��qa�lT0 k� ������2d q&�1D"3Q ��?    � ����m�_A�P ��1K��q|+� �ץ@�GHms��\gA��qa�lT0 k� ������2d q&�1D"3Q ��?    � ����m�_A�P ��1K��q|+� �ץ@�GHms��\gA��qa�lT0 k� ������2d q&�1D"3Q ��?    � ����m�_A�P ��1K��q|+� �ץ@�GHms��\gA��qa�lT0 k� �����2d q&�1D"3Q ��?    � ����n�_A�P ��2K��q|+� �ץ@�GHms��\gA��qa�lT0 k� �l �p 2d q&�1D"3Q ��?    � ����n�_A�P ��2K��q|+� �ץ@�GHmw��\gA��qa�lT0 k� �\�`2d q&�1D"3Q $�?    � ����n�_A�P ��2K��q|+� �ץ@�GHmw��\gA��qa�lT0 k� �`�d2d q&�1D"3Q ��?    � ����n�_K��P ��2K��q|+� �ץ@�GHmw��\gA��qa�lT0 k� �d�h2d q&�1D"3Q ��?    � ����o�_K��P ��2K��q|+� �ץ@�GHmw��\gA��qa�lT0 k� �h�l2d q&�1D"3Q ��?   � ����o.�_K��P ��2K��q|+� �ץ@�GHm{��\gA��qa�lT0 k� �l�p2d q&�1D"3Q ��?    � ����o.�_K��P ��2K��q|+� �ץ@�GHm{��\gA��qY�lT0 k� �p�t2d q&�1D"3Q ��?    � ��                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��>f ]�)�)� � � S;t   U @ 	   ���zp     SQ�����    ����             
 Z���         ��b     ��� 0		 
 
          c�   � �
	   ���zZ     b�����f    ���             :	 Z���         ���    ���    	!
           Oy�    	    ���     O�����Z    ���            	 Z��         �0     ���   H
           93   *      ��8G     9z���Y     )             	  Z��           � �     ���  0	 

          ]��  � �
	  .����     ]����B    ���	             Z	 Z��          ��    ���   @	
          ��S�  ��
     B�
i�    ��S��
i�                               ��              �  ���    8

 '            ���K          V�5�x    �����5�x                     Y  �� 
         (     ��B   0
&


          I2y        j��G     I2y��G                    	     �          
�     ��B   (
 
          �Ք         ~�m��    �Ք�m��       i            ���Z         0     ��J   0	
           i�/   9      � Uti     i�/ Uti                       �� O         	 �     ��@   H	$
          p��  H	     � ���     p�� ���                       
   O         
 .     ��@   03 
           ,��	      � �     , �                           
  �� L             a  ��@    P		 5                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          >�  ��        ����9  C� >?���t�  C����                    x                j  �       �                          >    ��       ���       >  ��           "                                                 �                         �����������
�5���m U � ������� 
 	               
   �  
 �"� ���C       %� `[� &d \� &� \� �$  g  �d g@ �� g`���J ����X ����J ����X � !d ] ��� ���� ����  ����. ����< ����J ����X � 
�\ W� �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �D �Q` � }`���� � ބ �`� � �^@ � _@  � �[� � \� � �j� � k� � �m@ � n@ �� �o� �� p� � �t� � u� �� w@ � �w` �$ x� �� �r@ �� s@���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �������� �� d  ������  
�fD
��L���"����D" � j  "  B   J jF�"      �j * , .��
��
��"   "D�j�
�� " �
� �  �  
�  O    ��     ���       O    ��     ���      ��    ��     ��m      ��  � ��   � � �         LL     �    ��        MM     �    ��        a�         �    ��  �"      ��0T ���        � �T ���        �        ��        �        ��        �   �     ��� ��        ��                          襩 4  
���                                     �                 ����             O�����%��   ����               18 Denis Savard ld                                                                                  2  1     �?cV �W c^ �k~ � k� � �K.O � K6W � K7G �K8G � 	K:O � 
K;R � �3 � �2 �K? �K/ �B�Q � B�a � B�I � B�L � B�R � B�T �B�E � B�U � B�M �kj4 � kr, �"�; � "�M ��7 �
�F �"�; � "�M � "�7 �!*�F*""� �* #"� �$� � 
� �m&*�.'"� �. ("�
)� � 
� 
� �,*� �-"� � ."�. �/� � 
�' �  "P q �  "J t �  "J v ~ 4"B y �  "J y �  "J { � 7"B | �  "J | �  "J | �  "K �@ ;"F �8<" �@ !� q8>" �@ !� q                                                                                                                                                                                                                         �� P         �     @ 
        �     _ P E a  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    �d~�f� ��������������������������������������������������������   �4, C   $ I� ��@(����n ��ł��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	        x    +      �   0$�J      ��                             ������������������������������������������������������                                                                                                                                 
       �    ���                      ��                  
   �������� ����������������������������������� ��������������� �� ������������ ������������������������������������ �� �� ��������� ������������� �� ������� ����  � ��������������������������������������� ���� ��� ����� � ������������                                       :    ��  D��J                                     ������������������������������������������������������                                                                       	                                                              	      �    ���                        �  �            
 	    �� ����� ��� ���� ��� ������������������������ � �� ������������ ������ ������������������ ����������� ������� � � ���������� ���������������� ������ ����������������������������������� �������� �����������������������������������                                                                                                                                                                                                                                                                                   	                                       �             


             �   }�                         ,�  HF                                   !6  Z                     �����������  	�  2�    ������������������������������������������������  �����  V��������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 8 F <                                  � �T� �\                                                                                                                                                                                                                                                                                       )n)n�  
                a      d      m      b      `            m                                                                                                                                                                                                                                                                                                                                                                                                               > �  >�  (�  (�  @  Bm'  ̆ F��d�k�����˶�c �V ����������������q�                ���D : � n          �   &  AG� �   �                    �                                                                                                                                                                                                                                                                                                                                        7 H          (             !��                                                                                                                                                                                                                            Y   �� �~ ���      �� \      �������� ����������������������������������� ��������������� �� ������������ ������������������������������������ �� �� ��������� ������������� �� ������� ����  � ��������������������������������������� ���� ��� ����� � �������������� ����� ��� ���� ��� ������������������������ � �� ������������ ������ ������������������ ����������� ������� � � ���������� ���������������� ������ ����������������������������������� �������� �����������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     @      @    �  >                       \     �   ����������      ��     T      �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �� ��  � ��     � ��   	 ��   p �� �� ��  � ��  � ��  �@ �� �� �z  �@���6 �$  �� ��   � ��   ��   ��     ��   � �� �� �    � �$ ^$  (   �   �� �� ��  �� �� �  �� �� �z � ��� �$ G �  ��G  �      �  ��   +�����������J  g���        f ^�         �� 2       +      ��>��������J���J��Q����      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                                         �� �����虙������(��������������񙙘�!                �  �������                           �       �  "(� """ �"" ""  "   �      �   �"��"""�"""�"""�"""�����������������������������������""�".�"/��"���!���.���/���-���""����������.���-������/�������   ��  �  .� /�� "�� "� "-�                                ""�  �(��""! ("" �"  �"   ����������������陙����.��� 陙/���.���"���"!��"��".���!♒""����������������̎���""�""",""/ �-� /� "�� "�� . /� �                    �                                           ""陂".��""� � �          �"(��(""������� ��        ""!�"!������������           ��     �                       wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  ""   "! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  ""   "! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!  " ! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        	�� ��� ��� ��� ��{ ��g �۶ �� ��  -�  �8 
3� D> 	D3 �C0˳ "+  ""  "   ��  �  ��  �  ��   ��  ��  wڐ kک g���w����ə�ͼ���܈��;��33̽�B��N�+0 ""@ B�  B$� K� ȋ  ʠ  +   "  �"" "�             �  �� �  ��  �   �� ��� ��       �                     �  �� �  �  �   �     ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                     ��� ���� ��    �     �                         � ���� ��   � � �           � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                              �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��                       "  .���"    �     �                       �   ��  ���  � �    �                                                                                                                                                     �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �                           � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ��л�� ���  �"  " ��"�""��"! � �  �   �   �   �                                                                                                                          �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                             �� ��������p��}` ��  �                        �   �   �                              ����������                                  "  .���"    �     �                         � ���� ��   � � �                                                                                                                                  "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��             �  �˰ ��� �wp ���                                                                                                                                                                �  ��� ��� ��Ъ�ݪ�	ڪ� ���	������������ �ۼ ��� 	�� �� �H�D��JE��E �� ���� ��� �� 	��+��+ـ"/ �"/ �  �    �            ��  �ː ̸� �ڋ ˽� ̻� ��� �̻ �˻�̻�����0���@��T3UUS3TK�8Dȸ�@�۰�ذ ً  ��  ��  )"� "" �"��� �� �            �   �   �   �   �                   �   ��     �               �  �� ���� ���  �    �       �  �  �  �  �  �   �                                     �   �           �   ̰  �˰                                                                                                                                                                                                                �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                            ��  ��  ��          ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ���     �     �                                                                                                                                                                                                  �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                    �   ��   ���  ��            �           �   �           "   "   "  �� ��                   ����������                                   � ��                  �  �˰ ��� �wp ���                                                                                                                                                                �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���          �     �  ��  ��   �                        �  ��            �   �    �                                ���� ��� ����                            ��  ��  ���                   ���                                                                                                                                                                                                    ��	����ɪ�ܙ����ݼ "-� "� J.��#��C>Z�C U�D �Z�#�U"�C"�� ���                �  �˰ ̻� �wp ׶� �vp �w� ɪ� ��� ��� �ۙ ��� �
� �" 0�" 0.�@ "�            ����˰ + �"  "" "  � �     �  �  ��  �   �               �   �   �   �   �   �   �@      �    �  �   �����������                   �   �                              �   �                      �������  ���    � ��  �   ��  �                  �       �                        �   ��  ���  � �    �                                                                                                                                       ̰ �� ̻ {�����vz� w��  ��  ��  ̘  	�  
� "��,̻�"�� "#3  34  D  
�  �  " "" """ ! ��  ��                               ˹� �ɩ ��� �͋ ��� ��� ��̀��Ȑ���лܹнȝ0ݙ�@43�PCD�@@E�@ E�@ U�� H�  K�  �   ��    �� "�" ���                          �  �   ��  �  ��                �   �   �   "   "   "  !�    ��                                 �   �                      �������  ���    �                    ��  ��  ���   �       �                        �   ��  ���  � �    �                               �   �                                                                                                    �  ��  ̽  ��  �w 
�� ���̹����	��̚���ȭ�̻������  ��  H� EU 4E C3  D;  ��  ��  ��  �  �  �   �  "  ��               �   �   �   �   ��  ��� ��� ��� ͻ���ة��ڌ�̽��˽����虚�DD��UT�"DUJ�3ET��DD��4M��ً�������۰��ـ+���+�ۿ��ۏ����"� �    �   �   �   ɀ  ��  ��         �    �  �       �                � ��� ��� ��  �                �   �     �   �           �  ��  ��  ��  ��� ��� ��� ��˰ɜ˰��˻�̻���������3���DDD�                                                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""��������D�M����""""�������D�M�M""""�����AMAD������""""��������D��""""������MM�����""""���������D�""""������������������""""������������������������"""$���4���4���4���4���4���4ffffffffffffffffff333DDDffffffffffffffffffffffff3333DDDDafaafffaffDDffff3333DDDDfFfFDfFFfFffdFffff3333DDDDfaffaffaffafffDfffff3333DDDDADAFaFadFfDffff3333DDDDafffDfdFdffff3333DDDDDDFFDfFFfdFffff3333DDDDAffAffaffafffDffffff3333DDDDffffffffffffffffffffffff3333DDDDfff4fff4fff4fff4fff4fff43334DDDD"""������������������""""������������������������""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""���������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��������������D�����3333DDDDI����D��DI����3333DDDDADAIA����D������3333DDDD��������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq?cV �W c^ �k~ � k� � �K.O � K6W � K7G �K8G � 	K:O � 
K;R � �3 � �2 �K? �K/ �B�Q � B�a � B�I � B�L � B�R � B�T �B�E � B�U � B�M �kj4 � kr, �"�; � "�M ��7 �
�F �"�; � "�M � "�7 �!*�F*""� �* #"� �$� � 
� �m&*�.'"� �. ("�
)� � 
� 
� �,*� �-"� � ."�. �/� � 
�' �  "P q �  "J t �  "J v ~ 4"B y �  "J y �  "J { � 7"B | �  "J | �  "J | �  "K �@ ;"F �8<" �@ !� q8>" �@ !� q3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������"��;�U�T��2�K�^�Z�G�R�R� � � � � � � � � ��=�@�����������������������������������������!��,�X�K�Z�Z��2�[�R�R� � � � � � � � � � ��=�@�����������������������������������������#��.�K�T�O�Y��<�G�\�G�X�J� � � � � � � � �=��;�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������=��;� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ������������������=�@� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������,�-��.�/�0�1�2������������������������� �!�"�3�4�#�#�#�#�#�#�#�#�$������������������%�&�'�(�)�)�)�)�)�)�)�)�)�)�*�+������������������5�6���7�8�9�:�;�<�=�>�?�������������������� �!�"�#�#�#�#�#�#�#�@�4�#�$������������������%�A�B�C�D�E�F�G�H�I�J�K�L�M�N�O�����������������P�Q�R�S�T�U�V�W�X�Y�W�Z�[�\�]�^��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            