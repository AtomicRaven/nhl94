GST@�                                                            \     �                                               2  �   8                  � 2���b�	 J���������������t���        >h      #    t���                                d8<n    �  ?     �����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    "�j��,  " ��
  �                                                                              ����������������������������������      ��    bb QQb  114 44c c   c      		 

       	   
       ��G �   ( (                 nhp ))1         888�����������������������������������������������������������������������������������������������������������������������������oo    gg                         ��                                                  ��            88 �����������������������������������������������������������������������������                                �j  j       R�   @  #   �   �                                                                                'w w  )n)h1p  ��    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    C�s�B9�8 q/�|/�E�P/�D@uE �����
���c��T0 k� �K��O�%�@2`QU8D"!  ��3    ��� {Dk�B8�4 q3�|/�E�H/��D8uE �����
���c��T0 k� �O��S�%�@2`QU8D"!  ��3    ��� |Dc�B8�0 q7�|/�E�D/�D0uE �����
���c��T0 k� �S��W�%�@2`QU8D"!  ��3    ��� }D[�B 7�, q?�|/�E�@/�D(uE �����R��c��T0 k� �[��_�%�@2`QU8D"!  ��3    ��� DS�A�6�( qC�|/�E�8/�DuE �����R��c��T0 k� �_��c�%�@2`QU8D"!  ��3    ��� �DC�A�5�  qO�|/�E�,/��DuB������R��c��T0 k� �k��o�%�@2`QU8D"!  ��3    ��� �D?�Q�4 qS�|/�D2(/��D uB������R��c��T0 k� �s��w�%�@2`QU8D"!  ��3    ��� �D7�Q�4 qW�|/�D2 0��D�uB������C�c��T0 k� �w��{�%�@2`QU8D"!  ��3    ��� �D/�Q�3 q_�|/�D20�߻I��uB������C�c��T0 k� �����%�@2`QU8D"!  ��3    ��� �D�Q�1 qg�|/�D21�߻I��uE ����C�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �D���0Q �o�|/�D21�߻I��uE ����C�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �D��/Q �s�|/�D22�߻I��uE {������c��T0 k� ����%�@2`QU8D"!  ��3    ��� �D��.Q �{�|/�D1�2�ۻI��uE ������c��T0 k� ����%�@2`QU8D"!  ��3    ��� �D��,P�
 ���|/�D1�3�׼I��uB��������c��T0 k� ����%�@2`QU8D"!  ��3    ��� �I���+P�	��|/�D1�4�ӼI��uB�������#�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �I����*P���|/�D1�4�ӼI��uB�������'�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �I����(P���|/�DA�5�ӼI��uB�������'�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �I����'P���|/�DA�5�ϼI��uB�������+�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �I���%P�A��|/�DA�7�˼I��uB�����/�c��T0 k� �ǈ�ˈ%�@2`QU8D"!  ��3    ��� �I��x#	��A��|/�DA�8�˼I��uB�����/�c��T0 k� �Ӈ�ׇ%�@2`QU8D"!  ��3    ��� �I��t"	��A��|/�E�8�˼I��uB�����3�c��T0 k� �߇��%�@2`QU8D"!  ��3    ��� �I��p 	��AË|/�E�9�˼I��uB�����3�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �I��h	��Aǋ|/�E�:�ǼI�xuB�����3�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �A��`	��A׌|/�E�<�ǼI�puB࣯��7�c��T0 k� ������%�@2`QU8D"!  ��3    ��� �A��\	��1ی|/�E�<�ǼI�luB࣭��7�c��T0 k� �����%�@2`QU8D"!  ��3    ��� �A��X	��1�|/�E�=�ǼI�huB৫��7�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �A��T	�� 1�|/�E�>üI�duB৩��7�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �A��P	�� 1�|/�E�?üI�`uB૧ b���7�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �A��L	�� 1�|/�E�x@ûI�\uB૥ b���7�c��T0 k� ����%�@2`QU8D"!  ��3    ��� �A���L	���!��|/�E�tAûI�XuB௣ b���7�c��T0 k� ���#�%�@2`QU8D"!  ��3    ��� �A���D	���"�|/�E�dD�ǺI�PuBೠ b���3�c��T0 k� �+��/�%�@2`QU8D"!  ��3    ��� �A���D	���"�|/�E�\E�˹I�LuBೞ ����3�c��T0 k� �/��3�%�@2`QU8D"!  ��3    ��� �E���@	���"�|/�E�XF�˹I�HuBො ����3�c��T0 k� �7��;�%�@2`QU8D"!  ��3    ��� �E����@	���B�|/�E�PG�˹I�HuBේ ����/�c��T0 k� �;��?�%�@2`QU8D"!  ��3    ��� �E����<		���B�|/�E�HH�˹I�DuE �� ����/�c��T0 k� �?��C�%�@2`QU8D"!  ��3    ��� �E����<	���B�|/�E�DJ�˹I�@uE �� ����/�c��T0 k� �G��K�%�@2`QU8D"!  ��3    ��� �E����<	���B#�|/�E�<K�ϸI�@uE ������+�c��T0 k� �K��O�%�@2`QU8D"!  ��3    ��� �F���8	���B'�|/�E�8L�ϸI�<uE Ó���C+�c��T0 k� �[��_�%�@2`QU8D"!  �3    ��� �F��8	���R3�|/�F,O�ӷI�<uE ǐ���C'�c��T0 k� �w��{�%�@2`QU8D"! ��?    ��� �F��8	���R7�|/�F$Q�׷I�8uEˎ���C#�c��T0 k� ����%�@2`QU8D"! ��?    ��� �F��8 	���R;�|/�F R�׶I�8uEˌ���C�c��T0 k� ����%�@2`QU8D"! ��?    ��� �D���;�	���R?�|/�FT�׶I�4uEϋ���C�c��T0 k� ����%�@2`QU8D"! ��?    ��� �D���?�	���RG�|/�FU�۵I�4uEӉ�����c��T0 k� ����%�@2`QU8D"! ��?    ��� �D���?�	���bK�|/�FV�۵I�4uEׇ�����c��T0 k� �Ǥ�ˤ%�@2`QU8D"! ��?    ��� �D���?�	���bO�|/�FX�ߵI�4uEۆ£���c��T0 k� �ק�ۧ%�@2`QU8D"! ��?    ��� �D���?�	���bS�|/�FZ�ߴI�4uE߄���c��T0 k� ����%�@2`QU8D"! ��?    ��� �F��C�	���bW�|/�F[�ߴI�0uE����c��T0 k� ������%�@2`QU8D"! ��?    ��� �F#��C�	���b[�|/�F ]��I�0uE����c��T0 k� ����%�@2`QU8D"!	 ��?    ��� �F'��G����b_�|/�F �^��I�0uE����c��T0 k� ����%�@2`QU8D"!
 ��?    ��� �F+��G����bc�|/�E��`��I�0uE��җ���c��T0 k� �#��'�%�@2`QU8D"!
 ��?    ��� �F/��K����bg�|/�E��a��I�0uE��җ����c��T0 k� �3��7�%�@2`QU8D"! ��?    ��� �E�3��O����bk�|/�E��c��A�0uE���ғ��� c��T0 k� �C��G�%�@2`QU8D"! ��?    ��� �E�7��O����bo�|/�E��d��A�0uE���ҏ��� c��T0 k� �S��W�%�@2`QU8D"! ��?    ��� �E�;��S�@��bs�|/�E��f��A�0uE���ҏ���c��T0 k� �c��g�%�@2`QU8D"! ��?    ��� �E�C��W�@��bw�|/�E��g��A�0uD��ҋ���c��T0 k� �s��w�%�@2`QU8D"! ��?    ��� �E�G��[�@��b{�|/�B��h��A�0uD��⇰��c��T0 k� �����%�@2`QU8D"! ��?    ��� �EK��_�@��b�|/�B��j��BA0uD��⃰��c��T0 k� �����%�@2`QU8D"! ��?    ��� �EO��_�@��b��|/�B��k��BA0uD������"���T0 k� �����%�@2`QU8D"! ��?    ��� �EW��c�@��b��|/�B��l��BA0uD������"���T0 k� �����%�@2`QU8D"! ��?    ��� �E[��g� ��b��|/�B��n��BA0uE���{���"���T0 k� �����%�@2`QU8D"! ��?    ��� �E_��o� ��b��|/�B��o��BA0uE�#��w���"���T0 k� ������%�@2`QU8D"! ��?    ��� �E�g��s� ��b��|/�B��p��BA0uE�'��s���"���T0 k� ������%�@2`QU8D"! ��?    ��� �E�k��w� ��b��|/�B��r��@0uE�/��o���)���T0 k� ������%�@2`QU8D"! ��?    ��� �E�o��{� �����|/�B��s��@0uE�3��k���)���T0 k� �����%�@2`QU8D"! ��?    ��� �E�w��� `�����|/�B��t �@4uE�;��g���)���T0 k� ����%�@2`QU8D"! ��?    ��� �E�{���� `�����|/�B��u �@4uE�?��c���)���T0 k� ����%�@2`QU8D"! ��?    ��� �D��ы� `�����|/�B��v �@4uE�C��_���)���T0 k� �+��/�%�@2`QU8D"! ��?    ��� �DӇ�я� `�����|/�B��x �B�4uEqK��[���)���T0 k� �;��?�%�@2`QU8D"! ��?    ��� �DӋ�ї� `�����|/�B��y �B�8uEqO�rW���)���T0 k� �K��O�%�@2`QU8D"! ��?    ��� �Dӓ�ћ������|/�B��z b�B�8uEqS�rW�¨)���T0 k� �[��_�%�@2`QU8D"! ��?    ��� �Dӗ�џ������|/�B��{ b�B�8uEq[�rS�¤)���T0 k� �k��o�%�@2`QU8D"! ��?    ��� �I�ѧ�� ���|/�B��| b�B�<uEq_�rO� )���T0 k� �{���%�@2`QU8D"! ��?    ��� �I�ѫ�� ���|/�B��} b�B�@uEqc�rK�)���T0 k� � �� %�@2`QU8D"! ��?    ��� �I�ѳ�� �Û|/�B��~ b�B�@uEqg�rG�)���T0 k� ����%�@2`QU8D"! (�?    ��� �I������ǜ|/�B�� ��B�DuEqo�rC�)���T0 k� $���%�@2`QU8D"! ��?    ��� �I������˝|/�B�� ��B�HuEqs�rC�)���T0 k� $�	��	%�@2`QU8D"! ��?    ��� �J�������ϝ|/�B�� ��B�HuEqw�r?�)���T0 k� $���%�@2`QU8D"! ��?    ��� �J�������Ӟ|/�B��� ��B�LuD�{�r;�)���T0 k� $���%�@2`QU8D"! ��?    ��� �J�������ן|/�B�� ��B�PuD��r7���)���T0 k� $���%�@2`QU8D"! ��?    ��� �J�������۠|/�B�� ��B�TuD���r7���)���T0 k� $���%�@2`QU8D"! ��?    ��� �J�������ߠ|/�B�  ��B�XuD���r3��|)���T0 k� �|��%�@2`QU8D"! ��?    ��� �I������ߠ|/�B� ��B�\uD���r/��x)���T0 k� �x�|%�@2`QU8D"! ��?    ��� �I�ô������|/�B�~2�B�`uD���r/��t)���T0 k� �t�x%�@2`QU8D"! ��?    ��� I�ô������|/�B�~2�B�duD���r+�bp)���T0 k� �p"�t"%�@2`QU8D"! ��?    ��� I�Ǵ������|/�B�~2�B�huD���r'�bl)���T0 k� �l%�p%%�@2`QU8D"!
 ��?    ��� I�Ǵ�����|/�B�~2�B�luD���r'�bh)���T0 k� 4h(�l(%�@2`QU8D"!	 ��?    ��� J˴������|/�E�~2�B�tuD���r#�bd)���T0 k� 4d+�h+%�@2`QU8D"! ��?    ��� J˴������|/�E�}"�B�xuD���r�b`)���T0 k� 4`.�d.%�@2`QU8D"! ��?    ��� J˴������|/�E� }"��B�|uD���r�b\)���T0 k� 4\1�`1%�@2`QU8D"! ��?    ��� Jϴ/�����|/�E�(}"��B��uD���r�RT )���T0 k� 4T8�X8%�@2`QU8D"! ��?    ��� I�ϴ7������|/�E�,}"��B��uD�����RP )���T0 k� �P;�T;%�@2`QU8D"! ��?    ��� I�ϴ?������|/�E�0|"��B��uD�����RL c��T0 k� �L>�P>%�@2`QU8D"! ��?    ��� I�ϴG������|/�E�8|��B��uD�����RH c��T0 k� �HA�LA%�@2`QU8D"! ��?    ��� I�ӴO���	���|/�E�<|��B��uD�ð��RD d�T0 k� �DD�HD%�@2`QU8D"!  ��?    ��� JӴc���
���|/�E�H{�B��uD�˴���;�d�T0 k� �<J�@J%�@2`QU8D"!  ,�?    ��� JӴ�k������|/�E�L{�BѴuD�˶��7��T0 k� $8M�<M%�@2`QU8D"!  ��?    ��� JӴ�s������|/�E�T{�BѸuD�Ϸ��/��T0 k� $4P�8P%�@2`QU8D"! ��?    ��� JӴ�{������|/�E�Xz�B��uD�ӹ��+��T0 k� $0T�4T%�@2`QU8D"! ��_    ��� JӴ���� ���|/�E�\z�B��uD�׻��#��T0 k� $,W�0W%�@2`QU8D"! ��_    ��� @cӴ�������|/�I1dz�B��uD�۽�R��T0 k� $(Z�,Z%�@2`QU8D"! ��_    �  @cӴ�������|/�I1ly��B��uD�����R���T0 k� � `�$`%�@2`QU8D"! ��_    �  @cӴ�������|/�I1py��B��uD��� ��R���T0 k� �c� c%�@2`QU8D"! ��_    �  @cӴ�������|/�I1ty��B��uD��� ��R���T0 k� �f�f%�@2`QU8D"! ��_    � 
 @cӴ���� ���|/�IAxy�#�B��uD��� ��Q����T0 k� �i�i%�@2`QU8D"! ��_    �  @�Ӵ����(���|/�IA|y�'�B��uD��� ��A����T0 k� �l�l%�@2`QU8D"! ��_    �  @�Ӵ����,��|/�IA�y�+�B�uD��� ��A����T0 k� Do�o%�@2`QU8D"! ��_    �  @�Ӵ����4��|/�IA�y�/�B�uD��� a��A����T0 k� Dr�r%�@2`QU8D"! ��_    �  @�Ӵ����8��|/�IA�y�3�B�uD��� a��A�����T0 k� Du�u%�@2`QU8D"! ��_    �  @�Ӵ����D��|/�I1�y�;�B�(uD��� a��A�����T0 k� D |�|%�@2`QU8D"! ��_    �  @�Ӵ����L��|/�I1�y�C�B�0uD��� a��A�����T0 k� ��� %�@2`QU8D"! )�_    �  �AӴ����P��|/�I1�y�G�B�<uD�����A�����T0 k� ����%�@2`QU8D"! ��_    �  �AӴ���T��|/�I1�y�K�B�DuD�����A�����T0 k� ����%�@2`QU8D"! ��_    �  �AӴ���\��|/�I1�y�O�B�LuD�����A�����T0 k� �����%�@2`QU8D"! ��_    �  �AӴ���`�߿|/�IA�y�S�B�TuD���������T0 k� �؀�܀%�@2`QU8D"! ��_    �  �C�ϴ���l"���|/�IA�y�_�B�huD���������T0 k� �Ȁ�̀%�@2`QU8D"! ��_    �   �C�ϳ��Ap#���|/�IA�y�c�B�puD���������T0 k� #���ā%�@2`QU8D"! ��_    � ! �C�ϳ�#�Ax%���|/�IA�y�k�B�|uD���������T0 k� #�����%�@2`QU8D"! ��_    � " �C�ϳ�+�A|&���|/�I1�y�o�B��uD���������T0 k� #�����%�@2`QU8D"! ��_    � # �C�˲�7�A�)���|/�I1�y�{�B��uD���������T0 k� #�����%�@2`QU8D"!  ��_    � $ �C�ǲ�?�A�+��|/�I1�y���B��uD���������T0 k� ������%�@2`QU8D"!  ��_    � % �C�Ǳ�C�A�,��|/�I1�ys��B��uD���������T0 k� ������%�@2`QU8D"!  -�_    � & �C�Ǳ�G�A�.��|/�IA�ys��B��uD�#��������T0 k� ������%�@2`QU8D"!  ��_    � ' �C�ð�S�A�1��|/�IA�ys��B��uD�'���{����T0 k� �p��t�%�@2`QU8D"!  ��_    � ( �C����W�A�3��|/�IA�ys��E�uD�+�B�s���T0 k� 3h��l�%�@2`QU8D"!  ��_    � ) �C����[�A�4��|/�IA�ys��E�vD�+�B�o���T0 k� 3`��d�%�@2`QU8D"!  ��_    � * �C����c�Q�6��|/�I1�ys��E�vD�/�B�k���T0 k� 3X��\�%�@2`QU8D"!  ��_    � + �C����k�Q�9��|/�I1�ys��E�vD�3�B�c���T0 k� 3H��L�%�@2`QU8D"!  ��_    � , �C����o�Q�;��|/�I1�ys��E��vD�7�B�_���T0 k� �@��D�%�@2`QU8D"!  ��_    � - �C����o�Q�<��|/�I1�ys��E�vD�4 B�W���	T0 k� �8��<�%�@2`QU8D"!  ��_    � . �C����w���@w�|/�@��ysǾE�uD�8B#�O���T0 k� �(��,�%�@2`QU8D"!  ��W    � / �C����{���ABo�|/�@��yc˽E�uD�<B#�AK���T0 k� �0��4�%�@2`QU8D"!  ��W    � 0 �C�������CBk�|/�@��ycӼBC(uD�<B#�AG���T0 k� �<��@�%�@2`QU8D"!  ��W    � 1 �C�������DBc�|/�@��yc׻BC0uEr@
B'�AC���T0 k� �D��H�%�@2`QU8D"!  ��W    � 2 �C���Ã���HBW�|/�@��yc߹BC@tErD"'�A7���T0 k� �X��\�%�@2`QU8D"!  ��W    � 3 �C���Ç���I�O�|/�A�yc�BCHtErD"+�A3���T0 k� �`��d�%�@2`QU8D"!  ��W    � 4 �C���Ç���K�G�|/�A�yc�BCPtErH"+�A/���T0 k� �h��l�%�@2`QU8D"!  ��W    � 5 �C���Ë���M�?�|/�A�yc�BCXsErH"/�A'���T0 k� �p��t�%�@2`QU8D"!  ��W    � 6 �C���Ï���P�3�|/�A�yc�BChsErL"3�A���T0 k� ������%�@2`QU8D"!  ��W    � 7 �C���ӏ���R�+�|/�A�yc�BCpsErL"7�A���T0 k� ������%�@2`QU8D"!  ��W    � 8 �CË�ӏ���T�#�|/�AQ�yc�BCxrErP"7�1���T0 k� ������%�@2`QU8D"!  ��W    � 9 �CË�ӏ���V��|/�AQ�yc��BC�rErP";�1���T0 k� ������%�@2`QU8D"!  ��W    � : �CÇ�ӓ���Y��|/�AQ�yc��BC�rErT""?�1���T0 k� ������%�@2`QU8D"!  ��W    � ; �CÇ�ӓ�� [��|/�AQ�yS��BC�rErX$�C�0����T0 k� ����%�@2`QU8D"!  ��W    � < �CÇ���� ]���|/�C�yS��BC�qEbX&�G�0����T0 k� ����%�@2`QU8D"!  ��W    � < �CÃ����_���|/�C�yS��BC�qEbX(�K�0����T0 k� ����%�@2`QU8D"!  ��W    � < �CÃ����a���|/�C�yS��BC�qEb\*�K�0� ��T0 k� ����%�@2`QU8D"!  ��W    � < �CÃ����e���|/�C�y��BC�qEb\.�S�0���T0 k� ��~��~%�@2`QU8D"!  ��W    � < �@������g���|/�C�y��BC�pEb\0�W�0���T0 k� ��~��~%�@2`QU8D"!  ��W    � < �@������i���|/�C�y��BC�pEb\2�[�0���T0 k� ��~��~%�@2`QU8D"!  �W    � < �@���C� BkA��|/�C�y��BC�pEb`4 b_�0���T0 k� ��~��~%�@2`QU8D"!  �W    � < �@��C�BnA��|/�C�yT�BC�pEb`8 bg�0�� T0 k� ��}��}%�@2`QU8D"!  ��W    � < �@��C�BpA��|/�C�yT�BC�oEb`: bk�0�� T0 k� ��}� }%�@2`QU8D"!  ��W    � < �@��C|BrA��|/�C�yT�BC�oEb`< bk�0�� T0 k� � }�}%�@2`QU8D"!  ��W    � < �@��C|BtA��|/�C�yT�BC�oEb`> bo�0�� T0 k� �}�}%�@2`QU8D"!  ��W    � < �@��CxBvA��|/�C�yT�BC�oEb`@ bs�0�	� T0 k� �|�|%�@2`QU8D"!  ��W    � < �@��Ct	BvA��|/�C�yT�BC�oEbdA bw�0�
�T0 k� �{�{%�@2`QU8D"!  ��W    � < �@��Ct
BuA��|/�C�yT�BD oEbdC b{� ���T0 k� �{�{%�@2`QU8D"!  ��W    � < �A�Cp2uA{�|/�C�yT�BDnA�dE b� ���T0 k� �z� z%�@2`QU8D"!  ��W    � < �A�Cl2tAs�|/�C�yT�BDnA�dG b� ���T0 k� � y�$y%�@2`QU8D"!  ��W    � < �A�3h2tAk�|/�C�|yT�BDnA�dI b�� ���T0 k� �$y�(y%�@2`QU8D"!  ��W    � < �A�3d2s1[�|/�C�tyT�BDnA�dL b�� ���T0 k� �,x�0x%�@2`QU8D"!  ��W    � < �AS�3`2s1S�!�/�DpyT�BD mA�dN b�� ���T0 k� �4x�8x%�@2`QU8D"!  ��W    � < �AS�3\ �s1K�!�/�DlyT�BD$lA�dO b�� ���T0 k� �8x�<x%�@2`QU8D"!  ��W    � < �AS��\ �s1C�!�/�DhyT�BD(kA�hQ b�� ���T0 k� �<w�@w%�@2`QU8D"!  ��W    � < �AS��X �s1;�!�/�D`yT�BD(jA�hS b�� ���T0 k� �@v�Dv%�@2`QU8D"!  ��W    � < �AS��T �r�3�!�/�D\yT�BD,iA�hT b�� ���T0 k� �Du�Hu%�@2`QU8D"!  ��W    � < �A���T �r�/�!�/�DXyT�BD0hA�hV b�� ���T0 k� �Dt�Ht%�@2`QU8D"!  ��W    � < �A���P br�'�!�/�DPyT�BD4gA�hW b�� ���T0 k� �Hs�Ls%�@2`QU8D"!  ��W    � < �A���L br��!�/�DLyT�BD4fA�hY b�� �|�T0 k� �Lr�Pr%�@2`QU8D"!  ��W    � < �A���L br��!�/�DHyT�BD8eA�hZ b�� �|�T0 k� �Lq�Pq%�@2`QU8D"!  ��W   � < �A���H  br��!�/�D@yT�BD<dA�h\ b�� �x�T0 k� �Pp�Tp%�@2`QU8D"!  ��W    � < �D���D" br��!�/�D<yT�BD<dA�h] b�� �t�T0 k� �To�Xo%�@2`QU8D"!  ��W    � < �D���D#�r��|/�I�4yT�BD@cA�l^ b�� �p�T0 k� �Xn�\n%�@2`QU8D"!  ��'    � < �D���@$�r���|/�I�0yT�BDDbA�l` b�� �l�T0 k� �Xm�\m%�@2`QU8D"!  ��'    � < �D���<&�r���|/�I�,yT�BDDaA�la b�� �l�T0 k� �\m�`m%�@2`QU8D"!  ��'    � < �D���<'� r���|/�I�(yT�BDH`A�lc b�� �h�T0 k� �`l�dl%�@2`QU8D"!  ��'    � < �D���8(� r���|/�I� yT�BDL_A�ld b�� �d�T0 k� �`k�dk%�@2`QU8D"!  ��'    � < �D���8*� r���|/�I�yT�BDL_A�le b�� �`�T0 k� �dj�hj%�@2`QU8D"!  ��'    � < �D���4+ $r���|/�I�yT�BDP^A�lf b�� �\�T0 k� �di�hi%�@2`QU8D"!  ��'    � < �D���4, $r���|/�I�yT�BDT]A�lh b�� �\�T0 k� �hi�li%�@2`QU8D"!  ��'    � < �D���0- $r�� |/�I�yT�BDT\A�li b�� �X�T0 k� �lh�ph%�@2`QU8D"!  ��'   � < �D���0/ $r��|/�I�yT�BDX\A�lj b�� �T�T0 k� �lg�pg%�@2`QU8D"!  ��'   � < �D���,0 $r��|/�I�yT�BDX[A�lk b�� �T�T0 k� �pf�tf%�@2`QU8D"!  ��'    � < �D���(1 (r��!�/�I�yT�BD\ZA�lm b�� �P�T0 k� �pe�te%�@2`QU8D"!  ��'    � < �D���(2 (rм!�/�I�yT�BD`ZA�pn b�� �L�T0 k� �te�xe%�@2`QU8D"!  ��'    � < �D���$3 (rи!�/�I� yT�BD`YA�po b�� �L�T0 k� �td�xd%�@2`QU8D"!  ��'    � < �D���$4 (rа!�/�I� yS��BD`XA�pp b�� �H�T0 k� �tc�xc%�@2`QU8D"!  ��'    � < �D��� 5 ,rЬ!�/�I��yS��BD`WA�pq b�� �D�T0 k� �tb�xb%�@2`QU8D"!  ��'    � < �D��� 6 ,rШ!�/�I��yS��BDdVA�pr b�� �D�T0 k� �xa�|a%�@2`QU8D"!  ��'    � < �D���7 ,rФ!�/�I��yS��BDdUA�ps b�� �@�T0 k� �|`��`%�@2`QU8D"!  ��'    � < �D���8 ,rР!�/�I��yS��BDdTA�pt b�� �< �T0 k� �|_��_%�@2`QU8D"!  ��'    � < �D���: ,rИ!�/�I��yS��BDdTA�pu b�� �< �T0 k� �|_��_%�@2`QU8D"!  ��'    � < �D���; 0rД	!�/�I��yS��BDdSA�pv b�� �8!�T0 k� �|^��^%�@2`QU8D"!  ��'    � < �D���< 0r0�
!�/�I��yS��BDhRA�pw b�� �8!�T0 k� ��]��]%�@2`QU8D"!  ��'    � < �D���< 0r0�
|/�I��yS��BDhQA�px b�� �4"�T0 k� ��\��\%�@2`QU8D"!  ��'    � < �D���= 0r0�|/�I��yS��BDhPA�py b�� �4"�T0 k� ��[��[%�@2`QU8D"!  ��'    � < �D���> 0r0�|/�I��yS�BDhPA�pz b�� �0"�T0 k� ��[��[%�@2`QU8D"!  ��'    � < �D���? 0r0�|/�I��yS�BDhOA�t{ b�� �,#�T0 k� ��Z��Z%�@2`QU8D"!  ��'    � < �D���@ 4r ||/�I��yS�BDlNA�t| b�� �,#�T0 k� ��Y��Y%�@2`QU8D"!  ��'    � < �D���A 4r x|/�I��yS�BDlNA�t} b�� �($�T0 k� ��Y��Y%�@2`QU8D"!  ��'    � < �D���B 4r t|/�I��yS�BDlMA�t~ b�� �($�T0 k� ��Y��Y%�@2`QU8D"!  ��'    � < �D���C 4r p|/�I��yS�BDlLA�t b�  �$$�T0 k� ��X��X%�@2`QU8D"!  ��'    � < �D���D 4r l|/�I��yS�BDlKA�t b�  �$%�T0 k� ��W��W%�@2`QU8D"!  ��'    � < �D���E 8r h|/�A��yS�BDpKA�t b� � %�T0 k� ��W��W%�@2`QU8D"!  ��'    � < �D���E 8r d|/�A��yS�BDpJA�t~ b� � &�T0 k� ��V��V%�@2`QU8D"!  ��'    � < �D���F 8r d|/�A��yS�BDpIA�t~ b� �&�T0 k� ��U��U%�@2`QU8D"!  ��'    � < �D��� G 8r `|/�A��yS�BDpIA�t~ b� �&�T0 k� ��U��U%�@2`QU8D"!  ��'    � < �D��� H 8r `|/�A��yS�BDpHA�t~ b� �'�T0 k� ��T��T%�@2`QU8D"!  ��'    � < �D��� I 8r \|/�A��yS�BDpHA�t} b� �'�T0 k� ��S��S%�@2`QU8D"!  ��'    � < �D����I 8r\|/�A��yS�BDtGA�t} b� �'� T0 k� ��S��S%�@2`QU8D"!  ��'    � < �D����J <rX|/�A��yS�BDtFA�t} b� �(� T0 k� ��R��R%�@2`QU8D"!  ��'    � < �D����K <rX|/�A��yS�BDtFA�t} b� �(� T0 k� ��R��R%�@2`QU8D"!  ��'    � < �D����L <rX|/�A��yS�BDtEA�t| b� �(� T0 k� ��Q��Q%�@2`QU8D"!  ��'    � < �D����L <rX|/�B@�yS�BDtEA�x| b� �)� T0 k� ��P��P%�@2`QU8D"!  ��'    � < �D����M�<r�T|/�B@�yS�BDtDA�x| b� �)� T0 k� ��P��P%�@2`QU8D"!  ��'    � < �D����N�<r�T |/�B@�yS�BDtDA�x| b�	 �)� T0 k� ��O��O%�@2`QU8D"!  ��'    � < �D����O�<r�T!|/�B@�yS�BDxCA�x| b�	 �*� T0 k� ��O��O%�@2`QU8D"!  ��'    � < �D����O�@r�T"|/�B@�yS�BDxBA�x{ b�
 �*� T0 k� ��N��N%�@2`QU8D"!  ��'    � < �D����P�@r�T#|/�B��yS߉BDxBA�x{ b�
 �*� T0 k� ��N��N%�@2`QU8D"!  ��'    � < �D����Q�@r�X$|/�B��yS߉BDxAA�x{ b� �*� T0 k� ��M��M%�@2`QU8D"!  ��'    � < �D����Q�@r�X%|/�B��yS߉BDxAA�x{ c  �+� T0 k� ��M��M%�@2`QU8D"!  ��'    � < �D����R�@r�X&|/�B��yS߉BDx@A�x{ c  �+�  T0 k� ��L��L%�@2`QU8D"!  ��'    � < �D����R�@r�X'|/�B��yS߉BDx@A�xz c  � +�$ T0 k� ��L��L%�@2`QU8D"!  ��'    � < �D����S�@r�\(|/�B��ySۉBD|?A�xz c � ,�$ T0 k� ��K��K%�@2`QU8D"!  ��'    � < �D��2�T�@r�\)|/�B��ySۉBD|?A�xz c � ,�$ T0 k� ��K��K%�@2`QU8D"!  ��'    � < �D��2�T�@r�\*|/�B��ySۊBD|>A�xz c ��,�$ T0 k� ��J��J%�@2`QU8D"!  ��'    � < �D��2�U�@r�`+|/�B��ySۊBD|>A�xz c ��,�$ T0 k� ��J��J%�@2`QU8D"!  ��'    � < �D��2�V�@r�d,|/�B��ySۊBD|>A�xz c ��-�$ T0 k� ��I��I%�@2`QU8D"!  ��'    � < �D��2�W�@r�d-|/�B��ySۊBD|=A�xz c ��-�$ T0 k� ��I��I%�@2`QU8D"!  ��'   � < �D��"�X�@r�h.|/�B� yS׊BD|=A�|y c ��-�$ T0 k� ��H��H%�@2`QU8D"!  ��'    � < �D��"�Y�@r�h.|/�B� yS׊BD|<A�|y c ��-�$ T0 k� ��H��H%�@2`QU8D"!  ��'    � < �D��"�Z�@r�l/|/�B�yS׊BD�<A�|y c ��.�$ T0 k� ��G��G%�@2`QU8D"!  ��'   � < �D��"�[�@r�p0|/�B�yS׊BD�;A�|y c ��.�$ T0 k� ��G��G%�@2`QU8D"!  ��'    � < �D��"�\�@r�t1|/�B�yS׊BD�;A�|y c ��.�$ T0 k� ��G��G%�@2`QU8D"!  ��'    � < �D��"�]�@r�x2|/�B�yS׊BD�;A�|y c ��.�$ T0 k� ��F��F%�@2`QU8D"!  ��'    � < �D��"�^�@r�|2|/�B�ySӊBD�:A�|y c ��/�$ T0 k� ��F��F%�@2`QU8D"!  ��'    � < �D��"�_�@r�|3|/�B�ySӊBD�:A�|y c ��/�$ T0 k� ��E��E%�@2`QU8D"!  ��'    � < �D��"�`�@r��4|/�B�ySӊBD�9A�|x c ��/�$!T0 k� ��E��E%�@2`QU8D"!  ��'    � < �D��"�a�@r��5|/�B�ySӋBD�9A�|x c ��/�$!T0 k� ��E��E%�@2`QU8D"!  ��'    � < �D���b�@q��5|/�B� ySӋBD�9A�|x c ��0�(!T0 k� ��D��D%�@2`QU8D"!  ��'    � < �D���c�@q��6|/�B�$ySӋBD�8A��x c ��0�(!T0 k� ��D��D%�@2`QU8D"!  ��'    � < �D�| �d�@q��7|/�B�(ySӋBD�8A��x c ��0�(!T0 k� ��D��D%�@2`QU8D"!  ��'   � < �D�|�e�@q��7|/�B�,ySϋBD�7A��x c ��0�(!T0 k� ��C��C%�@2`QU8D"!  ��'    � < �D�|�f�@q��8|/�B�0ySϋBD�7A��x c ��0�(!T0 k� ��C��C%�@2`QU8D"!  ��'    � < �D�|�g�@q��9|/�B�4ySϋBD�7A��x c ��1�(!T0 k� ��B��B%�@2`QU8D"!  ��'    � < �D�|�h�Dq��9|/�B�8ySϋBD|6A��x c ��1�(!T0 k� ��B��B%�@2`QU8D"!  ��'    � < �D�|	�i�Dq��:|/�B�@ySϋBD|6A��x c ��1�(!T0 k� ��B��B%�@2`QU8D"!  ��'    � < �D�|�j�Dqа;|/�B�DySϋBD|6A��w c ��1�(!T0 k� ��A��A%�@2`QU8D"!  ��'    � < �D�|�k�Dqи;|/�B�HySϋBD|5A��w c ��1�(!T0 k� ��A��A%�@2`QU8D"!  ��'    � < �D�| l�Dqм<|/�B�PySϋBDx5A��w c ��2�(!T0 k� ��A��A%�@2`QU8D"!  ��'    � < �D�|m�Dq��<|/�B�TySϋBDx5A��w c ��2�(!T0 k� ��@��@%�@2`QU8D"!  ��'    � < �D�|n�Dq��=|/�B�XySˋBDx5A��w c ��2�(!T0 k� ��@��@%�@2`QU8D"!  ��'    � < �D�|�o�Dq��>|/�B�`ySˋBDx4A��w c ��2�(!T0 k� ��@��@%�@2`QU8D"!  ��'    � < �D�|�o�Dq��>|/�B�dySˋBDx4A��w c  ��2�(!T0 k� ��@��@%�@2`QU8D"!  ��'    � < �LS|�p�Dq��?|/�B�lySˋBDt4A��w c  ��2�(!T0 k� ��?��?%�@2`QU8D"!  ��'    � < �LS|�q�Dq��?|/�B�pySˌBDt3A��w c  ��3�(!T0 k� ��?��?%�@2`QU8D"!  ��'    � < �LS|�q�Dq��@|/�B�xySˌBDt3A��w c  ��3�(!T0 k� ��?��?%�@2`QU8D"!  ��'    � < �LS|�r�Dq��@|/�B�|ySˌBDt3A��w c  ��3�(!T0 k� ��>��>%�@2`QU8D"!  ��'    � < �LS| � s�Dq��A|/�BфySˌBDt2A��v c  ��3�("T0 k� ��>��>%�@2`QU8D"!  ��'    � < �LS|"�(s�Dq��B|/�BьySˌBDp2A��v c$ ��3"("T0 k� ��>��>%�@2`QU8D"!  ��'    � < �LS|$�,t�Dq�B|/�BѐySǌBDp2A��v c$ ��3","T0 k� ��>��>%�@2`QU8D"!  ��'    � < �LS|%�0t�Dq�C|/�BјySǌBDp2A��v c$ ��4","T0 k� ��=��=%�@2`QU8D"!  ��'    � < �LS|'�4t�Dq�C|/�BѠySǌBDp1A��v c$ ��4","T0 k� ��=��=%�@2`QU8D"!  ��'    � < �LS|)�8u�Dq�D|/�B��ySǌBDp1A��v c$ ��4","T0 k� ��=��=%�@2`QU8D"!  ��'    � < �LS|*�<u�Dq� D|/�B��ySǌBDl1A��v c$ ��4","T0 k� ��<��<%�@2`QU8D"!  ��'    � < �LS|,�Du�Dq�(E|/�B��ySǌBDl1A��v c( ��4","T0 k� ��<��<%�@2`QU8D"!  ��'    � < �LS|.�Hu�Dq�,E|/�B��ySǌBDl0A��v c( ��4","T0 k� ��<��<%�@2`QU8D"!  ��'    � < �LS|/�Lu�Dq�4F|/�B��ySǌBDl0A��v c( ��4","T0 k� ��<��<%�@2`QU8D"!  ��'    � < �Lc|1�Pu�Dq�<F|/�B��ySǌBDl0A��v c( ��5","T0 k� ��;��;%�@2`QU8D"!  ��'    � < �Lc|2�Xu�Dq�@F|/�B��ySǌBDl0A��v c( ��5","T0 k� ��;��;%�@2`QU8D"!  ��'    � < �Lc|4�\u�Dq�HG|/�B��ySǌBDh/A��v c( ��5�,"T0 k� ��;��;%�@2`QU8D"!  ��'    � < �Lc|5�`u�Dp�LG|/�B��ySÌBDh/A��v c, ��5�,"T0 k� �|;��;%�@2`QU8D"!  ��'    � < �Lc|7�hu�Dp�TH|/�B��ySÌBDh/A��v c, ��5�,"T0 k� �|;��;%�@2`QU8D"!  ��'   � < �Lc|8�lu�Dp�XH|/�B��ySÌBDh/A��u c, ��5�,"T0 k� �|:��:%�@2`QU8D"!  ��'    � < �Lc|9�tu�Dp�`I|/�B��ySÌBDh/A��u c, ��5�,"T0 k� �|:��:%�@2`QU8D"!  ��'    � < �Lc|;�xu Hp�dI|/�K� ySÌBDh.A��u c, ��6�,"T0 k� �|:��:%�@2`QU8D"!  ��'    � < �Lc|<�|t Hp�lI|/�K�ySÍBDh.A��u c,  ��6�,"T0 k� �|:��:%�@2`QU8D"!  ��'    � < �Lc|>�t Hp�pJ|/�K�ySÍBDd.A��u c,  ��6�,"T0 k� �x:�|:%�@2`QU8D"!  ��'    � < �Lc|?�t Hp�xJ|/�K�ySÍBDd.A��u c,  ��6�,"T0 k� �x9�|9%�@2`QU8D"!  ��'    � < �Lc|@�s Hp�|K|/�K�ySÍBDd.A��u c0  ��6�,"T0 k� �x9�|9%�@2`QU8D"!  ��'    � < �Lc|A�s Hp��K|/�K�zSÍBDd-A��u c0! ��6�,"T0 k� �x9�|9%�@2`QU8D"!  ��'    � < �Lc|C�r�Ho��K|/�K�zSÍBDd-A��u c0! ��6"$,"T0 k� �x9�|9%�@2`QU8D"!  ��'    � < �Lc|D��r�Ho��L|/�K�zSÍBDd-A��u c0! ��6"$,"T0 k� �x9�|9%�@2`QU8D"!  ��'   � < �Lc|E��r�Ln��L|/�K� {SÍBDd-A��u c0! ��6"$,"T0 k� �x8�|8%�@2`QU8D"!  ��'    � < �Lc|F��q�Ln��L|/�K�${SÍBDd-A��u c0! ��7"$,"T0 k� �x8�|8%�@2`QU8D"!  ��'    � < �Lc|H��p�Lm��M|/�K�({SÍBD`,A��u c0" ��7"$,"T0 k� �t8�x8%�@2`QU8D"!  ��'    � < �Lc|I��p�Pm��M|/�K�,|S��BD`,A��u c0" ��7"$,"T0 k� �t8�x8%�@2`QU8D"!  ��'    � < �Lc|J��o�Pm��M|/�K�0|S��BD`,A��u c4" ��7"$,!T0 k� �t8�x8%�@2`QU8D"!  ��'    � < �Lc|K��n�Pl��N|/�K�4|S��BD`,A��u c4" ��7"$,!T0 k� �t8�x8%�@2`QU8D"!  ��'    � < �Lc|Ls�n�Tl��N|/�K�8}S��BD`,A��u c4" ��7"$,!T0 k� �t7�x7%�@2`QU8D"!  ��'    � < �Lc|Ms�m�Tk��N|/�K�<}S��BD`,A��u c4# ��7"$,!T0 k� �t7�x7%�@2`QU8D"!  ��'    � < �Lc|Ns�l�Tk��O|/�K�@}S��BD`,A��u c4# ��7"$,!T0 k� �t7�x7%�@2`QU8D"!  ��'    � < �Lc|Ps�j�Xj��O|/�K�H~S��BD`,A��u c4# ��7�,!T0 k� �t7�x7%�@2`QU8D"!  ��'    � < �Lc|QS�j�Xj��P|/�K�H~S��BD`+A��u c4# ��8�,!T0 k� �t7�x7%�@2`QU8D"!  ��'    � < �Lc|RS�i�Xj��P|/�K�L~S��BD`+A��u c4# ��8�,!T0 k� �t7�x7%�@2`QU8D"!  ��'    � < �Lc|SS�h�\i��P|/�K�PS��BD`+A��u c4$ ��8�,!T0 k� �t7�x7%�@2`QU8D"!  ��'   � < �Lc|TT g�\i��Q|/�K�TS��BD`+A��u c8$ ��8�,!T0 k� �t7�x7%�@2`QU8D"!  ��'    � < �Lc|UTf�\i��Q|/�K�XS��BD`+A��u c8$ ��8�,!T0 k� �t7�x7%�@2`QU8D"!  ��'    � < �Lc|VTf�`h��Q|/�K�\�S��BD`+A��u c8$ ��8�,!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �Lc|WTe�`h��R|/�K�\S��BD`+A��u c8$ ��8�,!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �Lc|XTd�`h��R|/�K�`S��BD`+A��u c8$ ��8�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �Lc|YTc�`g��R|/�K�dS��BD`+A��u c8% ��8�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �Lc|ZT$c�dg��R|/�K�dS��BD`+A��u c8% ��8�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �Lc|[T(b�dg�S|/�K�d~S��BD`+A��u c8% ��8�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �Lc|\T,a�df�S|/�K�d~S��BD`*A��u c8% ��9�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �Lc|]T4`�df�S|/�K�d~S��BD`*A��t c8% ��9�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �Lc|^T8`�hf�S|/�K�h~S��BD`*A��t c8% ��9�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �Lc|^d<_�he� T|/�K�h~S��BD`*A��t c<% ��9�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �LS|_d@^�he�(T|/�K�l~S��BD`*A��t c<& ��9�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �LS|`dH^�he�0T|/�K�l~S��BD`*A��t c<& ��9�(!T0 k� �t6�x6%�@2`QU8D"!  ��'    � < �LS|adL]�le�8T|/�K�l~S��BD`*A��t c<& ��9�(!T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �LS|bdP\�ld�@U|/�K�p~S��BD`*A��s c<& ��9�(!T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �LS|bdT\�ld�HU|/�K�p~S��BD`*A��s c<& ��9�(!T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �LS|cdX[�ld�PU|/�K�t~S��BD`*A��s c<& ��9�(!T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �D�|dd\[�ld�TU|/�K�t~S��BD`*A��s c<& ��9�( T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �D�|ed`Z�pe�\U|/�K�t~S��BD`*A��s c<' ��9�( T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �D�|fddY�te�dT|/�K�x~S��BD`*A��s c<' ��9�( T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �D�|gdhY�te�lT|/�K�x~S��BD`)A��r c<' ��:�( T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �D�|hdpX�xf�tT|/�K�|~S��BD`)A��r c<' ��:�( T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �E�|idtX�xf�xT|/�K�|~S��BD`)A��r c<' ��:�$ T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �E�|jdxW�|fS|/�K�|~S��BD`)A��r c@' ��:�$ T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �E�|kd|W�|gS|/�K��~S��BD\)A��r c@' ��:�$ T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �E�ld�V��gS|/�K��~S��BD\)A��r c@' ��:�$ T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �E�md�U��gҘS|/�K��~S��BD\)A��r c@' ��:�$ T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �F�nd�U��gҠR|/�K��~S��BD\)A��q c@( ��:�$ T0 k� �t5�x5%�@2`QU8D"!  ��'    � < �F�od�T��gҨR|/�K��~S��BD\)A��q c@( ��:�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �F�pd�T��gҰR|/�K��~S��BD\)A��q c@( ��:�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �F�rd�S��gҸR|/�K��~S��BD\)A��q c@( ��:�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �F�sd�R��g��R|/�K��~S��BD\)A��q c@( ��:�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �F�td�R��g��Q|/�K��~S��BD\)A��q c@( ��:�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��ud�Q��g��Q|/�K��~S��BD\)A��q c@( ��:�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��vd�P��g��Q|/�K��~S��BD\)A��q c@( ��:�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��xd�O��h��Q|/�K��~S��BD\)A��q c@( ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��yd�O��h��Q|/�K��~S��BD\)A��q c@) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��zd�N��h��P|/�K��~S��BD\)A��q c@) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��{d�M��h��P|/�B��~S��BD\(A��q c@) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��|d�M��h�P|/�B��~S��BD\(A��q cD) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��}d�L��h�P|/�B��~S��BD\(A��q cD) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��~d�K��h�P|/�B��~S��BD\(A��q cD) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��d�J��h� O|/�B��~S��BD\(A��q cD) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E���d�J��i�(O|/�B��~S��BD\(A��q cD) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E���d�I �i�0O|/�B��~S��BD\(A��q cD) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E���d�I �i�8O|/�B��~S��BD\(A��q cD) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��d�H �i�DO|/�K��}S��BD\(A��q cD) ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��d�G �i�LO|/�K��}S��BD\(A��q cD* ��;�$ T0 k� �t4�x4%�@2`QU8D"!  ��'    � < �E��d�G �i�TN|/�K��}S��BD\(A��q cD* ��;�$ T0 k� �t3�x3%�@2`QU8D"!  ��'    � < �E��~d�F �i�\N|/�K��}S��BD\(A��q cD* ��;�$ T0 k� �t3�x3%�@2`QU8D"!  ��'    � < �E��~d�F �i�dN|/�K��~S��BD\(A��q cD* ��;�$ T0 k� �t3�x3%�@2`QU8D"!  ��'    � < �E��}T�E �i�lN|/�K��~S��BD\(A��q cD* ��;�$ T0 k� �t3�x3%�@2`QU8D"!  ��'    � < �Cc�Ro��(���|/�F�le¯�B��9Ebg�3��Cc� �;T0 k� DO��S�%�@2`QU8D"! ��_    �  Cg�Ro��8���|/�F�pc¿�B��:Ebc�3���_� �:T0 k� $K��O�%�@2`QU8D"! ��_    �  Ck�Ro��@���|/�F�pb�ǧB��:Ebc�3���_� �:T0 k� $G��K�%�@2`QU8D"! ��_    �  Co�Ro��H���|/�@dpa�ӧB��:Eb_�3���_� �9T0 k� $C��G�%�@2`QU8D"! ��_    �  Cs�Ro��Pa��|/�@dp`�ۧB��:Eb_�����_� �8T0 k� $?��C�%�@2`QU8D"! ��_    �  Cw�Rl �Xa��|/�@dp_��B��;Eb[�����_� �8T0 k� $;��?�%�@2`QU8D"!  ��_    �  C{�Rl�da��|/�@dp]��B��;EbW�����[� �6T0 k� 43��7�%�@2`QU8D"!  ,�_    ��� C�Rl�la��|/�E�p\���E��<D2W�����[� �5T0 k� 4/��3�%�@2`QU8D"!  ��_    ��� C��Rl�ta��|/�E�p[��E��<D2S�����[� �4T0 k� 4+��/�%�@2`QU8D"!  ��_    ��� C��bl�|a��|/�E�pZ��E��<D2O�����W� �3T0 k� 4'��+�%�@2`QU8D"!  ��_    ��� C��bl��a��|/�E�pY��E��=D2O�����W� �2T0 k� 4#��'�%�@2`QU8D"! ��_    ��� C��bl	��1��|/�E�lV�'�E�>I�K�����S� �/T0 k� $���%�@2`QU8D"! ��_    ��� C#��bl��1��|/�E�lU%/�E�>I�K�����S���.T0 k� $���%�@2`QU8D"! ��_    ��� C#��bl��1��|/�E�lT%7�D�?I�G�����L ��,T0 k� $���%�@2`QU8D"! ��_    ��� C#��bl��1��|/�E�lR%?�D� ?I�G�����H��+T0 k� $���%�@2`QU8D"! ��_    ��� C#��bl��1��|/�E�lQ%G�D�,@I�G�����H��)T0 k� $���%�@2`QU8D"! ��_    ��� C#��bl��!��|/�E�lP%O�D�4@I�C�����D��(T0 k� D���%�@2`QU8D"! ��_    ��� I3��bl��#��|/�E�lM%_�E�DAI�C�ÿ��@��$T0 k� D���%�@2`QU8D"! ��_    ��� I3��rl��$��|/�E�lK%g�E�LBI�C�ӿ��<	��"T0 k� C����%�@2`QU8D"! (�    ��� �I3��rl��%��|/�E�lJ%o�E�XCI�?�ӻ��8�� T0 k� C����%�@2`QU8D"! ��    ��� �I3��rl��(��|/�E�hG%{�E�hDEb?�Ӵ �0��T0 k� �߀��%�@2`QU8D"!  ��    ��� �E���rl��)�{�|/�E�hE%��E�pEEb?�Ӱ �,��T0 k� �Ӏ�׀%�@2`QU8D"!  ��    ��� �E�ãrl��+�s�|/�E�hD%��E�xEEb?�Ӭ�(��T0 k� �ˀ�π%�@2`QU8D"!  -�    ��� �E�Ǣrl ��,�o�|/�E�dB%��E��FEb?�Ӭ�$��T0 k� ӿ��À%�@2`QU8D"!  ��    ��� �E�Ϣrl$��/�g�|/�E�`?%��Es�GEb?�Ӥ���T0 k� ���%�@2`QU8D"!  ��    ��� �B�ס	Rl&��0�c�|/�E�`=%��Es�HEb?�Ӡ���T0 k� ���%�@2`QU8D"!  ��    ��� �B�ۡ	Rl(��2�_�|/�E�\<%��Es�IEb?�Ӝ���T0 k� ���%�@2`QU8D"! ��    ��� �B��	Rl+��5�W�|/�E�X8%��Es�KEb?�Ӑ���T0 k� ��%�@2`QU8D"! ��    ��� �B��	Rl-��6�S�|/�E�X7%��Es�LEb?�ӌ���T0 k� �w~�{~%�@2`QU8D"! ��    ��� �B��	Rl/��7�O�|/�E�T5%��Es�MEb?��� ��
T0 k� �k~�o~%�@2`QU8D"! ��    ��� �B��	bl0��9�K�!�/�E�P4%��Es�NEb?������	T0 k� �_~�c~%�@2`QU8D"! ��    ��� �B���	bl3� ;�C�!�/�E�L1%çEs�QA�?��t	����T0 k� �K~�O~%�@2`QU8D"! ��    ��� �B��	bl4� =�C�!�/�E�H/%ǦEs�RA�?��p
����T0 k� �C~�G~%�@2`QU8D"! ��    ��� �B��	bl6� >�?�!�/�E�D.%#˦Es�SA�;��h
�� ��T0 k� �7}�;}%�@2`QU8D"! ��    ��� �B��	Rl7�?�;�!�/�E�@,%#ϦEs�UA�;��d�� �� T0 k� �+~�/~%�@2`QU8D"! ��    ��� �B��	Rl:�B�3�!�/�E�8)%#ۥEd XER;��X��"���T0 k� �~�~%�@2`QU8D"!  ��    ��� �B��	Rl;�C�/�!�/�E�4(%#ߤEdYER;��P��"���T0 k� �~�~%�@2`QU8D"!  ��    ��� �B��	Rl<�D�+�!�/�E�0&%#�EdZER7��L��"���T0 k� �~�~%�@2`QU8D"!  ��    ��� �B�'�	bl>�G�'�!�/�E�$$%#�Ed]ER3��<��#���T0 k� ��~��~%�@2`QU8D"!  ��    ��� �B�+�	bl?�H�#�|/�E� "%#�Ed _ER3��8�$c��T0 k� ��~��~%�@2`QU8D"!  /�    ��� �B�/�	bl@�I��|/�E�!%#�Ed$aER/��0�$c��T0 k� ��~��~%�@2`QU8D"!  ��    ��� �B�3�	blA� J��|/�E� %��Ed,bER/��(�$c��T0 k� ��~��~%�@2`QU8D"!  ��    ��� �B�;�	RlB� L�|/�E�%��Ed4eC�'���$c��T0 k� �~��~%�@2`QU8D"!  ��    ��� �B�?�	RlC��L�|/�E�%�Ed8gC�'���$c��T0 k� �~��~%�@2`QU8D"!  ��    ��� �B�C�	RlD��M�|/�E�%�Ed<iC�#���$c��T0 k� �~��~%�@2`QU8D"!  ��    ��� �B�G�	RlE��N�|/�E��%�Ed@jC����$c��T0 k� �~��~%�@2`QU8D"!  ��    ��� �B�O�	blF��O�|/�E��%�ETHnC�����$c��T0 k� �~��~%�@2`QU8D"!  ��    ��� �B�O�	blG��P�|/�E��%�ETLoC�����$c��T0 k� �~��~%�@2`QU8D"!  ��    ��� �B�O�	blG��P��!�/�E��%�ETHpC�����#c��T0 k� �w~�{~%�@2`QU8D"!  ��    ��� �B�O�	blH��Q��!�/�E��%$�ETDpC����
�#c��T0 k� �k~�o~%�@2`QU8D"!  ��    ��� �B�O�	blH��Q��!�/�E��%$�ETDpC����
�#c��T0 k� �c~�g~%�@2`QU8D"!  ��?    ��� �B�O�	RlI��R��!�/�E��%$�C�@pC����	�#c��T0 k� �W~�[~%�@2`QU8D"!  ��?    ��� �B�O�	RlI��R��!�/�E��%$�C�<pC������"c��T0 k� �O~�S~%�@2`QU8D"!  ��?    ��� �B�O�	RlI��Rp��!�/�E��%$�C�8pC�����|"c��T0 k� �C~�G~%�@2`QU8D"!  ��?    ��� �B�O�	RlJ��Rp��!�/�D��%$�C�0pC������x!c��T0 k� �/~�3~%�@2`QU8D"!  ��?    ��� �B�S�	blJ��Rp��!�/�D��%$�C�,qC������t!c��T0 k� �'�+%�@2`QU8D"!  ��?    ��� �B�S�	blJ��Rp��!�/�D��%$�C�$qC�����t c��T0 k� ��%�@2`QU8D"!  ��?    ��� �B�S�	blJ��Rp��!�/�D��%#��C� qC�����t c��T0 k� ��%�@2`QU8D"!  ��?    ��� �B�S�	blJ��Rp��|/�D�� c��C�qC�����p c��T0 k� ��%�@2`QU8D"!  ��?    ��� �@�S�	blK��Rp��|/�Ec� c��C�qC�����pc��T0 k� ���%�@2`QU8D"!  ��?    ��� �@�S�	RlK��Rp��|/�Ec� c��C�qP�����pc��T0 k� ����%�@2`QU8D"!  ��?    ��� �@�S�	RlK��Qp��|/�Ec� c��C�qP������pc��T0 k� ����%�@2`QU8D"!  ��?    ��� �@�S�	RlK��Q`��|/�Ec����C� qP������pc��T0 k� ����%�@2`QU8D"!  ��?    ��� �AS�	RlK��P`�|/�Ec����C��qP������pc��T0 k� ����%�@2`QU8D"!  ��?    ��� �AS�lK��P`�|/�Ec����C��rP������pc��T0 k� ����%�@2`QU8D"!  ��?    ��� �AS�lK��O`�|/�D3����C��rP������pc��T0 k� ���%�@2`QU8D"!  ��?    ��� ~AO�lK��O`�|/�D3|���C��rP������pc��T0 k� ���%�@2`QU8D"!  ��?    ��� |AO�lK��N`�|/�D3t���C��rP���ҋ�
Bpc��T0 k� ���%�@2`QU8D"!  ��?    ��� zATO�lK��M`�|/�D3p���D�rP���҇�
Bpc��T0 k� ���%�@2`QU8D"!  ��?    ��� xATK�RlK��L��|/�D3h���D�rP���҇�
Bpc��T0 k� ���%�@2`QU8D"!  ��?    ��� uATK�RlK��L��|/�D3d��D�rP���҃�
Bpc��T0 k� ���%�@2`QU8D"!  ��?    ��� sATG�RlK��J��|/�D3X��D�rP�����"pc��T0 k� �w�{%�@2`QU8D"!  ��?    ��� pE�G�RlK��I��|/�D3P��D�rP����{�"pc��T0 k� �o�s%�@2`QU8D"!  ��?    ��� mE�C��lK��H��|/�D3H��D�rP����{�"pc��T0 k� �c�g%�@2`QU8D"!  ��?    ��� jE�C��lK��G �|/�D3D��D�rP���{�"pc��T0 k� �[�_%�@2`QU8D"!  ��?    ��� hE�?��lK��F ߓ|/�D3<��D�sP�{��w�"pc��T0 k� �O�S%�@2`QU8D"!  ��?    ��� eE�;��lK��E ߓ|/�DC8��D�sP�w��w�2pc��T0 k� �G�K%�@2`QU8D"!  ��?    ��� cE�;��lK��D ߓ|/�DC0�߮D�sP�s��w�2pc��T0 k� �?�C%�@2`QU8D"!  ��?    ��� aE�7��lK��C ߓ|/�DC(�ۮD�sEQk��s�2pc��T0 k� �3�7%�@2`QU8D"!  ��?    ��� aD43��lK��A ے|/�DC$�ׯD�sEQg��s�2pc��T0 k� �#��'�%�@2`QU8D"!  ��3    ��� aD43��lJa�@�ے|/�DC�ׯDxsEQc��s�2pc��T0 k� ����%�@2`QU8D"!  ��3    ��� aD4/��lJa�?�ے|/�DC�ӰDlsEQ_��s�Bpc��T0 k� ����%�@2`QU8D"!  ��3    ��� aD4+��lJa�>�ۑ|/�DCSϰDdsEQ[��s�Bpc��T0 k� ����%�@2`QU8D"!  ��3    ��� aET#��lIa�;�ۑ|/�DC SǱDTsEQO�s�Btc��T0 k� ����%�@2`QU8D"!  ��3    ��� aET��lIa�:@ߐ|/�DB� SñDLsEQK�s�Btc��T0 k� �����%�@2`QU8D"!  ��3    ��� bET��lIa�9@ߐ|/�DB�!S��D@sEQC�s�Btc��T0 k� �����%�@2`QU8D"!  ��3    ��� cET��lHa�7@ߏ|/�Eb�"S��D8sEA?�s�Rtc��T0 k� �����%�@2`QU8D"!  ��3    ��� dET��lHa�6@ߏ|/�Eb�#S��D0tEA7�s�Rxc��T0 k� �����%�@2`QU8D"!  ��3    ��� eET�blGa�5@ߎ|/�Eb�$S��C�$tEA3�s�Rxc��T0 k� �����%�@2`QU8D"!  ��3    ��� fET�blFQ�3@�|/�Eb�%㫳C�tEA/�s�Rxc��T0 k� ���%�@2`QU8D"!  ��3    ��� gC��blFQ�2P�|/�Eb�%㣳C�tEA'�s�R|
c��T0 k� ��~�~%�@2`QU8D"!  ��3    ��� hC���bhDQ�/P�|/�Eb�'㗴C� tEA��w�R�c��T0 k� ��|�|%�@2`QU8D"!  ��3    ��� iC���bhDQ�.P�|/�Eb�(㓴C��tEA��w�R�c��T0 k� �|�|%�@2`QU8D"!  ��3    ��� jC��bdCQ�-P�|/�Eb�)㏵C��tEA��{�R�c��T0 k� �{�{%�@2`QU8D"!  ��3    ��� kC��bdBQ�,��|/�Eb�*ㇵC��tEA��{�R�c��T0 k� ��%�@2`QU8D"!  ��3    ��� lC��2dAQ�*��|/�Eb�,ヶC��tEA���
Ҍc��T0 k� ����%�@2`QU8D"!  ��3    ��� mC�ߩ2`A�|)��|/�ER�-�{�C��tE0����
Ґc��T0 k� ����%�@2`QU8D"!  ��3    ��� nC�۩2`@�x(��|/�ER�.�s�C��tE0�����
Ґc��T0 k� ����%�@2`QU8D"!  ��3    ��� oC�Ϫ2\>�l&���|/�ER�0�g�C�tE0�����
Ҙc��T0 k� ����%�@2`QU8D"!  ��3    ��� pC�Ǫ2X=�h$���|/�ER�0�_�C�tE0��	��
Ҝc��T0 k� ����%�@2`QU8D"!  ��3    ��� qC�ê2T=�d#��|/�ER�0�[�C�tE0��	��
Ҡ c��T0 k� ����%�@2`QU8D"!  ��3    ��� rC�2L=�`"��|/�ER|0�S�C�uE0��	��
Ҥ c��T0 k� ���#�%�@2`QU8D"!  ��3    ��� sC�2H<�\!��|/�ERx0�K�C�uE0��	��
ҫ�c��T0 k� �#��'�%�@2`QU8D"!  ��3    ��� tC�2D<�X ��|/�ERp0�C�C�uE0��	��
ү�c��T0 k� �'��+�%�@2`QU8D"!  ��3    ��� uC�28;�P��|/�C�h/�3�C�xuE0��	��
һ�c��T0 k� �/��3�%�@2`QU8D"!  ��3    ��� vC�B4;�L��|/�C�d/�+�C�puE0��	"��
��c��T0 k� �3��7�%�@2`QU8D"!  ��3    ��� wC�B,;�H��|/�C�\/�#�C�huE0��	"��
���c��T0 k� �7��;�%�@2`QU8D"!  ��3    ��� xC�B(:�D�#�|/�C�X/��C�\uE ��	"��
���c��T0 k� �;��?�%�@2`QU8D"!  ��3    ��� yC�B :�@�'�|/�C�P/��C�TuE ��	"��
���c��T0 k� �C��G�%�@2`QU8D"!  ��3    ��� z                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \���8 ]�'�'� � 
�� }�  [ Z     � ��     ~N� ���    �z�             M Z �          �p�     ��� 0
% 	           E��   � �	    �#�     F�#��    �e��             Q Z �         ��    ��� 0
 
          i�Z            ��     i�� �y;    sI             
  Z �           �     ���   8          N�I   Z Z     ��g     N�� ٠�     !/            ( Z �          M��     ��� P
	
         ��-�  ��	      .��
    ��-���
                               ���                  ���    P              ~�  � �
     B �0�     ~� ��!     ��         # 	  Z �          ���     ���   8

          ���   U       V �@    ��2 ��     G��              b��          ��     ��@   (
          (l� $ $       j�`     (v��M    �o��                �        }P     ��H  8�           qy�        ~ ��"     q�� �v�    ��b            
��          ��     ��@   	@
           *]�         � Ѧ     *I� љ�    2 �                  �         	 �      ��@   H
$
          ;ϩ        ���r�     ;����~     ��X            
    A �         
 �     ��@   H!	           W� ��      �	�      [:	    ����                      ���u             �  ��@      0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          3��  ��        ���  �� 3���  ���o��                   x                j  �       �                          3    ��        �       3             "                                                �                          �# � �� � � � ���	�� 	           
     
  [   �� 8)�J       D� `[� Dd d  D� d  D� d@ � i@ � i` A$ _����. ����< ����J ����X ����X � �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0� ���� ����� � � }`���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���� �  <���  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    "�j�� , " �
� �  �  
�  (    ��     �       i��  ��     � �       (    ��     �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �'��      ��4T ���        � �T ���        �        ��        �        ��        �   *�    ��
}���        ��                         T�) ,  ���                                     �                 ���� 
           (���%��   < �                 16 Pat Verbeek son y   4:34                                                                        4  4     �&C&	KB5-KH;KL;k~*0 k�: �c� �
c� � �	C � 
C  � C! � C"  �	J�4 � J�< � J�4 � J�, � c� � �c� � � c� � �	� � �	� � �� � �� � �kj � � kr � � � � � � � �B� �B� �B� � � B� � B� � �!"� � � ""� � �#� � �$
� �J%"�J &"�/:'"�:(*�, �)"� � � *"� � �+� � �,
� � u-" � �." � u/" � }0!� � u1" � u2* � � 3*HT � 4*KD � 5)�T �6*\ � 7*OT �8*(\ �9**l �:*8d � ;*Gd � <*Et =*Pd>"|- *lR@�R 
�                                                                                                                                                                                                         �� R @      �    @ 
        �     ] P E b  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    ��   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, >  6 ��	 ��@d��@��A���d�	�~��������                                                                                                                                                                                                                                                                                                                   @�                                                                                                                                                                                                                                                    c  	  $    ��  D�J    	  F�  	                           ������������������������������������������������������                                                                       
                                                         	          �      �      �                �  �          	  
 	 
 	 	 ��������������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� �                         
           "    ��  H�J       �                             ������������������������������������������������������                                                                                                                                           �        �      �        �    ��              
 	  
	 
 	 	 ����� ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� �������������           x                                                                                                                                                                                                                                        
                                                                     �             


           �   }�                                                                   'u                     ��������������������  N�������������  N�����������������    ��������  N�  N������������������������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww N @ 0 
              	                  � '1՚ �\                                                                                                                                                                                                                                                                                    )n)h1p  ��                    c      m               W       m                               ��                                                                                                                                                                                                                                                                                                                                                                       � � �  � ��  � ��  � (��  � (��  EZm:  �N z����������$����������������D����������yy          :  ���? :�� 		        	 �   & AG� �   �   
           � �                                                                                                                                                                                                                                                                                                                                      p B C    �     p                !��                                                                                                                                                                                                                            Y   �� �� ����      �� B 	     ��������������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ������ ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� �������������   �� �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    4      /   �  3                       B     �   ���������J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p����  �( �    � �$      �f ��     �f �$ ^$ �@      ����� ��   �����    ����0 ��   ����0 �$ ^$       �   | 
s� �� | 
s� �$ ^$�� l � ��� �� � ��� [ �2   A��A  �      �      /�������2����  g���         f ^�         ��M <      /      �������2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                               s   D   O   w   w   v   u   f   T   �   �              3@  DDp ��4 ��tp��wpO�tpdfwGfeTwfeWwfUFwdUFweTfp�DDp���p���@�w�p   C   D   O   D   w   u   U   U  F  d  f   f   D   �   �   �DD ���7���uP��e`O�V ffg ffG Ufw UU� FUN dFw ffp DDp ��p ��@ w�p  C4 4D@O�C���O�Dt�GVfeVfdFfdFfdUfffUfffwFff�DDD���� ���                    0   G   W   W   U   E   E   w   �   �   @    fg D� O�� �� w�}�w��}����������M���M���M��������y�                    �   �   �   �   �   �   �   �   ~   w       ���w���w���~���~�DMw�������������y�                        w���w}��wt��wt��w}M�����������   M   M   ~�  p�  p   p   p      �   �   �   �               vd  eVp ffpw�Op���w���G���M�}�                                     v   ub  ub  f   `   P               "  f  U` wfP        p   p   p   p   p   p   p   p                               C4 �y�                              f  vU`vf`D�O������p}�w�  ?�  ?�  ?�  33  3#                                      f  Ug                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "! ""! " "" """ "!   " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               ""   "! " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "! ""! " "" """ "!   " ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                     �  �  ��  8�  5I  5U  3U  DT  EZ UJ T� �J� ����+�""""�""//��          ��wɪ�pɪ��ɪ��̙�н��н̽Ѝɚݣ��"�<̲�;���0"�0  ="  ""  "/  /�� ���  �����                               �� �� �� ���          �.���       �  �      �  ��  �  ��  �              �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                      "  .���"    �     �                                                                                                                                                                                    ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     �  �  �  ��  �  �  �  ��  �             �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   ��  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �   �   �                .  ���� �                           �     �                                                                                                                                                                                                 �  �  ��  8�  5I  5U  3U  DT  EZ UJ T� �J� ����+�""""�""//��          ��wɪ�pɪ��ɪ��̙�н��н̽Ѝɚݣ��"�<̲�;���0"�0  ="  ""  "/  /�� ���  �����                               �� �� �� ���          �.���       �  �      �  ��  �  ��  �            �  �   �   ��  �                                  �� �� ��               �  �  �     �   �  �  �                                    ��  ��  ���                                                                                                                                                                                                        �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                                        "  "(��ȩ�ܚ��ۊ����� ��  �   �   �   �   �� ��� ̻� ˽� ��� �w� �������������������������� �̻ ���         �   �       �   �   "" �+� Ȼ� ɫ� ɨ� ��                �� �I��3 ��D 
UD 
UD TD  T�  ˸  ��  �� ̰ �+ ��"/ �"/  ����  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �   �   �                .                      ��  ��  ���              �  �˰ ��� �wp ���                                                                                                                                                                                     �  ɪ� ɪ� ̚� �ȍ ͷ  "�  "� .( 3># �4�
�T��T�"�UN"�UN(�Dɜ� ʨ����, � /�������� � ��                                ��  ��  ��  g}  �א vz� gz� ̊� �ɩ 8̜ D<� T� @��  �� ɀ ��  ��  "   .          �  ��� �������  ��                           "  "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����        ��� �  ��     �                                    �  �� �                         ����     �   �  �  �  ��  �   �                                                                                                             �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   �   �"  ""  !� �� ��  �               �   ������  ��                   �                        ���� ��� ����          �   �   �   �  �  �  �  �           �  ��� ݼ� w{� �װ vw�    �   ��  ���  � �    �                                                                                                                                       �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��  ��  ��� ���                                                �   ���                            �   �                                                                                                                         	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                                   ��                     �   �                      �������  ���    �                    ��  ��  ���     ��   �  ��  �  �  �         � �������������  �                                �   �                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �        �  ��  ��  ww  ��  vv  w"   "   "  �� ��                   ����������                      �  ������� ��                        ���                                                                                                                                                                                           �  ��� ܽи�؀  � ˚ �̹�̹�˹�˻ܻ��ܘ��܉���D���U�D�J�N T�� D�  T�  �  ��  �� �� ,ث"���"��� ���۝� {�� ��  ��� ��(�������� ˸� ɀ  ��  ��� �̀ �̈ �� ���虎�(���"��� ��� � �/�����              �   �   �   �   �   ��                                          �� ��� ��� ��  �                         �   �                     �   ��� �̰         �   �  �  �   �               �   �                                                    �   �   �   �   �   �                                                                                                                                                �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��           	 
          
        ((((((( 
	(((( ����������������             ! " # $ % & '   ( $ % ) ! " # * ('(&(%($(#("(! (((���������������� + , -   . / 0 1  	 2         3       4 (((((((2	10/(.(-(,(+���������������� 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5����������������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<���������������� L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L����������������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq&C&	KB5.KH;KL;k~*0 k�: �c� �
c� � �	C � 
C  C! � C"  �J�< � J�< � J�4 � J�, � c� � �c� � � c� � �	� � �	� � �� � �� � �kj � � kr � � � � � � � �B� �B� �B� � � B� � B� � �!"� � � ""� � �#� � �$
� �J%"�J &"�/:'"�:(*�, �)"� � � *"� � �+� � �,
� � u-" � �." � u/" � }0!� � u1" � u2* � � 3*HT � 4*KD � 5)�T �6*\ � 7*OT �8*(\ �9**l �:*8d � ;*Gd � <*Et =*Pd>"|- *lR@�R 
�L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������ �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������#� ��9�K�Z�X��5�R�O�S�G� � � � � � � � � � �/�.�7�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.�����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������/�.�7� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� �� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�A�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                