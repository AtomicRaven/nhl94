GST@�                                                           �e�                                                      � �� N     �  ��  1         ����e ����J����������� �������        �g     #    ����                                d8<n    �  ?     h����  �
fD�
�L���"����D"��   " `  J  jF��    "�j "����
��
��     �j�� 
   ��
  4�                                                                              ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������=  0b  4  11                                         �  �  �  �                  $  
          = �����������������������������������������������������������������������������                                ��  �       ��   @  #   �   �                                                                                '       )n)n1n  
$    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE 9 �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �,AMS\L$,?�ttE���Y|,  �@� �� c4# �S��!T0 k� ������&�1D"3Q	E1 4#Q  ��   �  ��,AMS\L$,?�xtE��Y|,  �@� �� c4# �S��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��,AMS`L$0>�xtE��Y|,  �@� �� c4$ �S��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��,AMS`L$0>�|tE��Y|,  �@� �� c4% �S��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��,AMSdL$4=��tD��Y|,  �@� �� c8% �S��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��,AMSdL$4=��sD��Y|,  �@� �� c8& �S��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��,AMchL$8<��sD��Y|,  �@� �� c8' �W��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0AMchL$<;��sD�#�Y|,  �@� �� c8( �W��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0AMchL$<;��sE�'�Y|,  �@� �� c<( �W��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0AMclL$<;��sE�/�Y|,  �@� �� c<) �W��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMclL@:��sE�3�Y|,  �@� �� c<) �W��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMclL@:��sE�;�Y|,  �@� �� c<* �W��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMcpLD9��sE�?�Y|,  �@� �� c<* �W��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMcpLD9��sE�G�Y|,  �@� �� c@+ �W��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMSp LH8��sE�K�Y|,  �@� �� c@+ �[��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMSt LH8��sE�S�Y|,  �@� �� c@, �[��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMSt!C�H8��sB�W�Y|,  �@� �� c@, �[��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMSt"C�L7��sB�_�Y|,  �@� �� c@- �[��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMSx"C�L7��sB�g�Y|,  �@� �� cD- �[��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��0BMSx#C�L7��sB�h Y|,  �@� �� cD. �[��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BMSx$C�L6��sB�p Y|,  �@� �� cD. �[��!T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BMSx$E�L6��sLpxY|,  �@� �� cD/ �[��"T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BMS|%E�L5��sLp|Y|,  �@� �� cD/ �[��"T0 k� ������&�1D"3Q	E1 4#Q  ��   �  ��4BD�|&E�L5��sLp�Y|,  �@� �� cD0 �[��"T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BD�|&E�L5��sLp�Y|,  �@� �� cH0 �_��"T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BD��'E�L5��rLp�Y|,  �@� �� cH1 �_��"T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BD��(E�L5��rLp�Y|,  �@� �� cH1 �_��"T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BD��)E�L5��rLp�Y|,  �@� �� cH1 �_��"T0 k� ������&�1D"3Q	E1 4#Q  ��   �  ��4BEs�)E�H5��rLp�Y|,  �@� �� cH2 �_��"T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BEs�*E�H5��rLp�Y|,  �@� �� cH2 �_��"T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BEs�+E�H5��rLp�Y|,  �@� �� cH3 �_��"T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BEs�,D4D5��rLp�Y|,  �@� �� cH3 �_��"T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��4BEs�-D4D5��rLp�Y|,  �@� �� cH4 �_��"T0 k� �����&�1D"3Q	E1 4#Q  ��    �  ��4BEc�.D4@5��rLp�Y|,  �@� �� cH4 �_��"T0 k� �����&�1D"3Q	E1 4#Q  ��    �  ��4BEc�/D4@5��rLp�Y|,  �@� �� cH5 �_��"T0 k� �{���&�1D"3Q	E1 4#Q  ��   �  ��4BEc�0D4<6��rL��Y|,  �@� �� cH5 �_��"T0 k� �{���&�1D"3Q	E1 4#Q  ��    �  ��8BEc�1D4<6��rL��Y|,  �@� �� cD5 �c��"T0 k� �w��{�&�1D"3Q	E1 4#Q  ��    �  ��8BEc�2D486��rL��Y|,  �@� �� cD6 �c��"T0 k� �w��{�&�1D"3Q	E1 4#Q  ��    �  ��8BD3�4D447��rL��Y|,  �@� �� cD6 �c��"T0 k� �s��w�&�1D"3Q	E1 4#Q  ��    �  ��8BD3�5DD47��rL��Y|,  �@� �� cD7 �c��"T0 k� �s��w�&�1D"3Q	E1 4#Q  ��    �  ��8BD3�6DD07��rL��Y|,  �@� � cD7 �c��"T0 k� �o��s�&�1D"3Q	E1 4#Q  ��    �  ��8BD3�7DD,8��rL��Y|,  �@� � cD8 �c��"T0 k� �o��s�&�1D"3Q	E1 4#Q  ��    �  ��8BD3�9DD,9��rL��Y|,  �@� � cD8 �c��"T0 k� �k��o�&�1D"3Q	E1 4#Q  ��    �  ��8BD3�:DD(9��rL��Y|,  �@� � cD8 �c��"T0 k� �k��o�&�1D"3Q	E1 4#Q  ��   �  ��8BD3�;DD$:��rL��Y|,  �@� � cD9 �c��"T0 k� �g��k�&�1D"3Q	E1 4#Q  ��    �  ��8BD3�<DD :��rL��Y|,  �@� � cD9 �c��"T0 k� �g��k�&�1D"3Q	E1 4#Q  ��   �  ��8BDC�>DD;��rL��Y|,  �@� � cD: �c��"T0 k� �c��g�&�1D"3Q	E1 4#Q  ��    �  � 8BDC�?DD<��rL��Y|,  �@� � cD: �c��"T0 k� �c��g�&�1D"3Q	E1 4#Q  ��    �  � 8BDC�ADD<��rL��Y|,  �@� � cD: �c��"T0 k� �_��c�&�1D"3Q	E1 4#Q  ��    �  � 8BDC|BDD=��rL��Y|,  �@� � cD; �c��"T0 k� �[��_�&�1D"3Q	E1 4#Q  ��    �  � 8BDC|CDT>��rL��Y|,  �@� � cD; �g��"T0 k� �[��_�&�1D"3Q	E1 4#Q  ��    �  � 8BDC|EDT?� rL� Y|,  �@� � cD< �g��"T0 k� �W��[�&�1D"3Q	E1 4#Q  ��   �  � 8BDCxFDT@�rL�Y|,  �@� � c@< �g��"T0 k� �W��[�&�1D"3Q	E1 4#Q  ��    �  ��8BDCtHDT A�rL�Y|,  �@� � c@< �g��#T0 k� �S��W�&�1D"3Q	E1 4#Q  ��    �  ��8BDCtIDS�A�rL�Y|,  �@� � c@= �g��#T0 k� �S��W�&�1D"3Q	E1 4#Q  ��    �  ��<BDCpKDS�B�rL�Y|,  �@� � c@= �g��#T0 k� �O��S�&�1D"3Q	E1 4#Q  ��    �  ��<BDClMDS�C�rL�Y|,  �@� � c@= �g��#T0 k� �O��S�&�1D"3Q	E1 4#Q  ��    �  ��<BDSlNDS�D� rL�Y|,  �@� � c@> �g��#T0 k� �K��O�&�1D"3Q	E1 4#Q  ��    �  ��<CDShPDS�E�$rL�Y|,  �@� � c@> �g��#T0 k� �K��O�&�1D"3Q	E1 4#Q  ��    �  ��<CDSdRDS�G�,rL�Y|,  �@� � c@> �g��#T0 k� �G��K�&�1D"3Q	E1 4#Q  ��    �  ��<CDS`SDS�H�0rL�Y|,  �@� � c@? �g��#T0 k� �G��K�&�1D"3Q	E1 4#Q  ��    �  ��<CDS`UDc�I�8rL� Y|,  �@� � c@? �g��#T0 k� �C��G�&�1D"3Q	E1 4#Q  ��    �  ��<CEc\WDc�J�<rL�$Y|,  �@� � c@? �g��#T0 k� �C��G�&�1D"3Q	E1 4#Q  ��    �  ��<CEcXXDc�K�DqL�(Y|,  �@� � c@@ �g��#T0 k� �?��C�&�1D"3Q	E1 4#Q  ��    �  ��<CEcTZDc�L�HqL�(Y|,  �@� � c@@ �g��#T0 k� �?��C�&�1D"3Q	E1 4#Q  ��    �  ��<CEcP\Dc�M�PqL�,Y|,  �@� � c@@ �g��#T0 k� �;��?�&�1D"3Q	E1 4#Q  ��    �  ��<CEcL^ES�O�XqL�0Y|,  �@� � c@A �g��#T0 k� �;��?�&�1D"3Q	E1 4#Q  ��    �  ��<CEcH_ES�P�\qL�4Y|,  �@� � c@A �k��#T0 k� �7��;�&�1D"3Q	E1 4#Q  ��    �  ��<CEcDaES�Q�dqL�4Y|,  �@� � c@A �k��#T0 k� �7��;�&�1D"3Q	E1 4#Q  ��    �  ��<CEc@cES�R�lqL�8Y|,  �@� � c@A �k��#T0 k� �3��7�&�1D"3Q	E1 4#Q  ��    �  ��<CES<eES�S�tqL�<Y|,  �@� � c@B �k��#T0 k� �3��7�&�1D"3Q	E1 4#Q  ��    �  ��<CES4gES�T�xqL�<Y|,  �@� � c@B �k��#T0 k� �/��3�&�1D"3Q	E1 4#Q  ��    �  ��<CES0hES�U߀qL�@Y|,  �@� � c@B �k��#T0 k� �/��3�&�1D"3Q	E1 4#Q  ��    �  ��<CES,jES�W߈qL�DY|,  �@� � c@B �k��#T0 k� �+��/�&�1D"3Q	E1 4#Q  ��    �  ��<CES(lES�XߐqL�DY|,  �@� � c<C �k��#T0 k� �+��/�&�1D"3Q	E1 4#Q  ��    �  ��<CES mC�YߘqL�HY|,  �@� � c<C �k��#T0 k� �'��+�&�1D"3Q	E1 4#Q  ��    �  ��<CESoC�|ZߠqLqLY|,  �@� � c<C �k��#T0 k� �'��+�&�1D"3Q	E1 4#Q  ��    �  ��<CESqC�t[ߨqLqLY|,  �@� � c<C �k��#T0 k� �'��+�&�1D"3Q	E1 4#Q  ��    �  ��<CESrC�p\߰qLqPY|,  �@� � c<D �k��#T0 k� �#��'�&�1D"3Q	E1 4#Q  ��    �  ��<CEStC�h]߸qLqPY|,  �@� � c<D �k��#T0 k� �#��'�&�1D"3Q	E1 4#Q  ��    �  ��<CESuES`^��qLqTY|,  �@� � c<D �k��#T0 k� ���#�&�1D"3Q	E1 4#Q  ��    �  ��@CEB�wESX_��qLqXY|,  �@� � c<D �k��#T0 k� ���#�&�1D"3Q	E1 4#Q  ��    �  ��@CEB�xESP`��qD�XY|,  �@� � c<E �k��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CEB�yESH`��qD�\Y|,  �@� � c<E �k��#T0 k� ����&�1D"3Q	E1 4#Q  ��   �  ��@CEB�{ES@a��qD�\Y|,  �@� � c<E �k��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CEB�|ES8b��qD�`Y|,  �@� � c<E �k��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CEB�}EC,c��qD�`Y|,  �@� � c<F �k��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CEB�~EC$d��qLqdY|,  �@� � c<F �k��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CEB�ECe� qLqhY|,  �@� � c<F �k��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CEB̀ECe�qLqhY|,  �@� � c<F �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CEBĀECf�qLqlY|,  �@� � c<F �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CE2�ECf�qLqlY|,  �@� � c<G �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CE2�EB�g�$qLqpY|,  �@� � c<G �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CE2�EB�g�,qLqpY|,  �@� � c<G �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CE2�~EB�h�4qLqtY|,  �@� � c<G �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CE2�~EB�h�<qLqtY|,  �@� � c<G �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CE2�}EB�h�HqLqxY|,  �@� � c<H �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CE2�|E2�i�PqL�xY|,  �@� � c<H �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@CE2�|E2�i�XqL�|Y|,  �@� � c<H �o��#T0 k� ����&�1D"3Q	E1 4#Q  ��    �  �\�5@��A���\��A+�Z��\�A��-W���PW�"s��T0 k� �;��?�&�1D"3Q	E1 4#Q  ��    �����\�5@��A���\��A+�Y}�\�A��-W���PW�"s��T0 k� �G��K�&�1D"3Q	E1 4#Q  ��    �����\�5@��A���\��A'�Y}�\�A��-[�ǋPW�"s��T0 k� �S��W�&�1D"3Q	E1 4#Q  ��    �����\�5@��A���\��A'�Y}�\�A��-[�ˋPS�"s��T0 k� �c��g�&�1D"3Q	E1 4#Q  ��    �����\�5@�A��\��A'�Y}�\�A��-[�ϋPP 3��T0 k� �o��s�&�1D"3Q	E1 4#Q  ��    �����\�5@�A��\��A#�Y}#�\�A��-_�ӌPP 3��T0 k� �{���&�1D"3Q	E1 4#Q  ��    �����\�5@�A�{�\��A#�Y}'�\�A��-_�یPP 3��T0 k� ������&�1D"3Q	E1 4#Q  ��    �����\�5@�A�{�\��A#�Y}+�\�A��-c�ߌPP 3��T0 k� ������&�1D"3Q	E1 4#Q  ��    �����\�5@�A�w�\��A�Y}/�\�A��-c��PP 3��T0 k� ������&�1D"3Q	E1 4#Q  ��    �����\�5@�A�w�\��A�Y}7�\�A��.c��PL 3��T0 k� ������&�1D"3Q	E1 4#Q  ��    �����\�5@�A�w�\��A�Y};�\�A��.g��PL 3��T0 k� ������&�1D"3Q	E1 4#Q  ��    �����\�5@�A�s�\��A�Y}?�\�A��.g��PL 3��T0 k� �˃�σ&�1D"3Q	E1 4#Q  ��    �����\�5@�A�s�\��A�Y}C�\�A��.g��PL 3��T0 k� �׃�ۃ&�1D"3Q	E1 4#Q  ��    ��� \�5@�A�o�\��A�Y}G�\�A��.k���PL 3��T0 k� ����&�1D"3Q	E1 4#Q  ��    ��� \�5@�A�o�\��A�Y}O�\�A��.k���PL 3��T0 k� ����&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�o�\��A�Y}S�\�A��.k���PH 3��T0 k� ������&�1D"3Q	E1 4#Q  ��    ��� 
\�6@�A�k�\��A�Y}W�\�A��.o���PH 3��T0 k� ����&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�k�\��A�Y}[�\�A��.o���PH 3��T0 k� ����&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�g�\��A�Y}_�\�A��.o���PH 3��T0 k� �#��'�&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�g�\��A�Y}c�[��A��.s���PH 3��T0 k� �/��3�&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�g�\��A�Y}g�[��A��.s���PH 3��T0 k� �;��?�&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�c�\��A�Y}k�[��A��.s���PH 3��T0 k� �O��S�&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�c�\��A�Y}o�[��A��.w��#�PD 3��T0 k� �W��[�&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�c�\��A�Y}s�[��A��.w��'�PD 3��T0 k� �[��_�&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�_�\��A�Y}w�[��A��.w��3�PD 3��T0 k� �_��c�&�1D"3Q	E1 4#Q  ��    ��� \�6@�A�_�\��A�Y}{�[��A��.{��?�PD 3��T0 k� �_��c�&�1D"3Q	E1 4#Q  ��    ��� \�6E�A�_�\��A�Y}�[��A��.{��G�PD 3��T0 k� �S��W�&�1D"3Q	E1 4#Q  ��    ��� \�6E�A�[�\��A�Y}��[��A��.{��S�PD 3��T0 k� �K��O�&�1D"3Q	E1 4#Q  ��    ��� \�6E�A�[�\��A�Y}��[��A��.{��_�PD 3��T0 k� �G��K�&�1D"3Q	E1 4#Q  ��    ��� \�6E#�A�[�\��A�Y}��[�A��.��k�PD 3��T0 k� �C��G�&�1D"3Q	E1 4#Q  ��    ��� \�6E#�A�W�\��A�Y}��[�A��.��k�P@ 3��T0 k� �C��G�&�1D"3Q	E1 4#Q  ��    ��� \�6FO'�A�W�\��A�Y}��[�A��.�w�P@ 3��T0 k� �G��K�&�1D"3Q	E1 4#Q  ��    ��� \�6FO'�A�W�\��A�Y}��[�A��.���P@ 3��T0 k� �K��O�&�1D"3Q	E1 4#Q  ��    ��� \�6FO+�A�S�\��A�Y}��[�A��.����P@ 3��T0 k� �O��S�&�1D"3Q	E1 4#Q  ��    ��� \�6FO+�A�S�\��A�Y}��[�A��.����P@ 3��T0 k� �S��W�&�1D"3Q	E1 4#Q  ��    ��� \�6FO/�A�S�\��A��Y}��[�A��.����P@3��T0 k� �S��W�&�1D"3Q	E1 4#Q  ��    ��� \�6FO/�A�O�\��A��Y}��[�A��.����P@3��T0 k� �W��[�&�1D"3Q	E1 4#Q  ��    ��� \�6F?3�A�O�\��A��Y}��[�A��/����P@3��T0 k� �W��[�&�1D"3Q	E1 4#Q  ��    ��� \�6F?3�A�O�\��A��Y}��[�A��/����P@3��T0 k� �[��_�&�1D"3Q	E1 4#Q  ��    ��� \�6F?7�A�O�\��A��Y}��[�A��/����P@3��T0 k� �[��_�&�1D"3Q	E1 4#Q  ��    ��� \�6F?7�A�K�\��A��Y}��[�A��/��ǔP<3��T0 k� �_��c�&�1D"3Q	E1 4#Q  ��    ��� \�6F?;�A�K�\��A��Y}��[�A��/��ϔP<3��T0 k� �k��o�&�1D"3Q	E1 4#Q �    ��� \�6F_;�A�K�\��A��Y}��[�A��/��וP<3��T0 k� �s��w�&�1D"3Q	E1 4#Q ��    ��� \�6F_?�A�K�\��A��Y}��[�A��/��ߕP<3��T0 k� �����&�1D"3Q	E1 4#Q ��    ��� \�6F_?�A�G�\��A��Y}��[�A��/���P<3��T0 k� ������&�1D"3Q	E1 4#Q ��    ��� \�6F_C�A�G�\��A��Y}Ã[�A��/���P<3��T0 k� ������&�1D"3Q	E1 4#Q ��    ��� #\�6F_C�A�G�\��A��Y}ǃ[�A��/����P<3��T0 k� ������&�1D"3Q	E1 4#Q	 ��    ��� '\�6FoG�A�G�\��A��Y}˃[�A��/����P<3��T0 k� ������&�1D"3Q	E1 4#Q
 ��    ��� +\�6FoG�A�C�\��A��Y}˃[�A��/���P<3��T0 k� ������&�1D"3Q	E1 4#Q ��    ��� /\�6FoG�A�C�\��A��Y}τ[�A��/���P<3��T0 k� �ã�ǣ&�1D"3Q	E1 4#Q ��    ��� 2\�6FoK�A�C�\��A��Y}ӄ[߫A��/���P<3��T0 k� �Ϧ�Ӧ&�1D"3Q	E1 4#Q ��    ��� 5\�6FoK�A�C�\��A��Y}ׄ[߫A��/���P83��T0 k� �ۨ�ߨ&�1D"3Q	E1 4#Q ��    ��� 8\�7FoO�A�?�\��A��Y}ׄ[߫A��/���P83��T0 k� ����&�1D"3Q	E1 4#Q ��    ��� ;\�7FoO�A�?�\��A��Y}ۄ[߫A��/��'�P83��T0 k� �����&�1D"3Q	E1 4#Q ��    ��� >\�7FoO�A�?�\��A��Y}߅[߫A��/��/�P83��T0 k� �����&�1D"3Q	E1 4#Q ��    ��� A\�7FoS�A�?�\��A��Y}߅[۫A��/��3�P83��T0 k� ����&�1D"3Q	E1 4#Q ��    ��� D\�7FoS�A�?�\��A��Y}�[۫A��/��;�P83��T0 k� ����&�1D"3Q	E1 4#Q ��    ��� G\�7FoS�A�;�\��A��Y}�[۫A��/���G�P83��T0 k� ���#�&�1D"3Q	E1 4#Q ��    ��� J\�7FoW�A�;�\��A��Y}�[۫A��/���S�P83��T0 k� �+��/�&�1D"3Q	E1 4#Q ��    ��� M\�7FoW�A�;�\��A��Y}�[۫A��/���_�P83��T0 k� �7��;�&�1D"3Q	E1 4#Q ��    ��� P\�7FoW�A�;�\��A��Y}�[׫A��/���o�P83��T0 k� �C��G�&�1D"3Q	E1 4#Q ��    ��� S\�7Fo[�A�;�\��A��Y}�[׫A��/���{�P83��T0 k� �O��S�&�1D"3Q	E1 4#Q ��    ��� V\�7Fo[�A�7�\��A��Y}�[׫A��/�����P83��T0 k� �W��[�&�1D"3Q	E1 4#Q ��    ��� Y\�7Fo_�A�7�\�A��Y}��[׫A��/�����P83��T0 k� �c��g�&�1D"3Q	E1 4#Q ��    ��� \���A���@���k�@�Y�  ��@�����]�����3� T0 k� �˺�Ϻ&�1D"3Q	E1 4#Q ��/    ����n���A���@���k�@�Y�  ��@�����]�����3� T0 k� �˺�Ϻ&�1D"3Q	E1 4#Q  /�/    ����l���A���@���k�@�Y�  ��@�����]�����3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����j���A���B����k�@�Y�� ��@����]�����3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����h���A���B����k�@�Y�� ��@����������3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����f���A���B����k�@�Y�� ��@����������3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����d���A���B����k�@�Y�� ��@����������3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����b���A���B����k�@�Y�� ��@����������3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����`L��BL��B���Lk�BL�Y����A���������3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����^L��BL��B���Lk�BL�Y����A���������3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����\L��BL��B�úLk�BL�Y����A���������3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����ZL��BL��B�úLk�BL�Y����A���������3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����XL��BL��B�ǺLk�BL�Y����A���������3� T0 k� ������&�1D"3Q	E1 4#Q ��/    ����V ��Dܧ�O˺�k�D��Y����A\�������M��3� T0 k� ������&�1D"3Q	E1 4#Q  ��/    ����T ��Dܧ�O˺�k�D��Y����A\����M��M��3� T0 k� ������&�1D"3Q	E1 4#Q  ��/    ����S ��Dܧ�O˺�k�D��Y����A\����M��M��3� T0 k� �����&�1D"3Q	E1 4#Q  ��/    ����R ��Dܧ�OϺ�k�D��Y����A\����M��M��3� T0 k� �{���&�1D"3Q	E1 4#Q  ��/    ����Q ��Dܧ�OϺ�k�D��Y����A\����M��M��3� T0 k� �w��{�&�1D"3Q	E1 4#Q  ��/    ����P l��Dܧ�OӺ�k�P��Y����A�����M��M��3� T0 k� �o��s�&�1D"3Q	E1 4#Q  /�/    ����N l��Dܧ�O׺�k�P��Y����A�������� ��3� T0 k� �k��o�&�1D"3Q	E1 4#Q  ��/    ����M l��Dܧ�O׺�k�P��Y����A�������� ��3� T0 k� �g��k�&�1D"3Q	E1 4#Q  ��/    ����L l��D짌Oۺ�k�P��Y����A����#���� ��3� T0 k� �_��c�&�1D"3Q	E1 4#Q  ��/    ����JL��D짍Oߺ�k�Q�Y����D����#���� ��3� T0 k� �[��_�&�1D"3Q	E1 4#Q  ��/    ����IL��D짎O��k�Q�Y����D����#�������3� T0 k� �O��S�&�1D"3Q	E1 4#Q  ��D    ����HL��D짎O��k�Q�Y����D����#�������3� T0 k� �G��K�&�1D"3Q	E1 4#Q  ��D    ����GL��D짏O��k�Q�Y����D����#������3� T0 k� �C��G�&�1D"3Q	E1 4#Q  ��D    ����F,��F��O��k�Q�Y����D����#������3� T0 k� �?��C�&�1D"3Q	E1 4#Q  ��D    ����E,��F��O��k�P��Y����D����#������3� T0 k� �;��?�&�1D"3Q	E1 4#Q  ��D    ����D,��F��O��k�P��Y����D����#������3� T0 k� �7��;�&�1D"3Q	E1 4#Q  ��D    ����D,��F��O��k�P��Y����D����#������3� T0 k� �3��7�&�1D"3Q	E1 4#Q  ��D    ����D,��F��O��o�P��Y����D����#������3� T0 k� �3��7�&�1D"3Q	E1 4#Q  ��D    ����D,��E���O��o�B\�Y���ߜD����#������3� T0 k� �3��7�&�1D"3Q	E1 4#Q  ��D    ����D,��E���O��o�B\�Y���ߝD����#������3� T0 k� �3��7�&�1D"3Q	E1 4#Q  ��D    ����D,��E���O��o�B\�Y���ߟD����������3� T0 k� �3��7�&�1D"3Q	E1 4#Q  ��D    ����D,��E���O���o�B\�Y���ۢD������ǩ�#�3� T0 k� �7��;�&�1D"3Q	E1 4#Q  ��D    ����D���E���B����o�B\�Y���ۣD������˩�'�3� T0 k� �7��;�&�1D"3Q	E1 4#Q  ��D    ����D���E���B����s�B\�Y���ץD������ϩ�+�3� T0 k� �7��;�&�1D"3Q	E1 4#Q  ��D    ����D���E���B���{�B\�Y���ӨD�����ש�3�3� T0 k� �;��?�&�1D"3Q	E1 4#Q  ��D    ����D���E���B���{�B\#�Y���ӪEm����۩�7�3� T0 k� �;��?�&�1D"3Q	E1 4#Q  ��D    ����D���E���B����B\'�Y���ϫEm������;�3� T0 k� �?��C�&�1D"3Q	E1 4#Q  ��D    ����D���E���B��܃�B\'�Y���ϭEm������?�3� T0 k� �C��G�&�1D"3Q	E1 4#Q  ��D    ����E���E���B��܋�Bl/�Y���ǰEm�����K�3� T0 k� �G��K�&�1D"3Q	E1 4#Q  ��D    ����F���E���B��܏�Bl/�Y��|ǲEm������O�3� T0 k� �K��O�&�1D"3Q	E1 4#Q  ��D    ����G���B���B��ܓ�Bl3�Y��|ôEm������W�3� T0 k� �O��S�&�1D"3Q	E1 4#Q  ��D    ����H���B���B��ܗ�Bl7�Y��|��Em�����[�3� T0 k� �O��S�&�1D"3Q	E1 4#Q  ��D    ����I,��B�ÛB�'�ܣ�Bl?�Y��|��Em
�����g�3� T0 k� �W��[�&�1D"3Q	E1 4#Q  ��D    ����J,��B�ǛB�+����Bl?�Y��|��D=�����k�3� T0 k� �[��_�&�1D"3Q	E1 4#Q  ��D    ����K,��E˛B�3����BlC�Y�����D=�����s�3� T0 k� �_��c�&�1D"3Q	E1 4#Q  ��D    ����L,��EϛB�7����BlG�Y�����D=���#��{�3� T0 k� �c��g�&�1D"3Q	E1 4#Q  ��D    ����M,�EלB�C����BlO�Y�����D=���3�އ�3� T0 k� �k��o�&�1D"3Q	E1 4#Q  ��D    ����N,�EߜB�G����B|S�Y�����E����;�ދ�3� T0 k� <w��{�&�1D"3Q	E1 4#Q �D    ����S,�E�B�O����B|W�Y�����E����?�ޓ�3� T0 k� <�����&�1D"3Q	E1 4#Q ��O    ����X,�E�B�[����B|_�Y�����E����O�ޣ�3� T0 k� <�����&�1D"3Q	E1 4#Q ��O    ����],�B��B�c����B|c�Y�����E����W�ާ�3� T0 k� <�����&�1D"3Q	E1 4#Q ��O    ����b 	B���B�g����H�g�Y��|��E����_�ޯ�3� T0 k� ������&�1D"3Q	E1 4#Q	 ��O    ����g
B���B�o�	��H�g�Y��|��E�!���g�޷�3� T0 k� ������&�1D"3Q	E1 4#Q ��O    ����lB��B��	��H�g�Y��|��E�&���w�	��3� T0 k� ������&�1D"3Q	E1 4#Q ��O    ����qB��B̓�	��H�k�Y��|��E}(����	��3� T0 k� ������&�1D"3Q	E1 4#Q ��O    ����vB��B͋�	��H�k�Y��	|��E}*�����	��3� T0 k� ������&�1D"3Q	E1 4#Q ��O    ����z B��B͓�	�H�k�Y��	|��E},�����	��3� T0 k� ����&�1D"3Q	E1 4#Q ��O    ����~(B�+�Bͣ�	-�H�k�Y�#�	|��E}1�����	��3� T0 k� ���#�&�1D"3Q	E1 4#Q ��O    �����0B�3�Bͫ�	-�H�o�Y�#�	|��E}3������	.��3� T0 k� �+��/�&�1D"3Q	E1 4#Q ��O    �����8B�7�Bݳ�	-�Io�Y�#�	|��E}6������	.��3� T0 k� M7��;�&�1D"3Q	E1 4#Q ��O    �����<B�?�Bݻ�	-�Io�Y�#�	���E}8������	.��3� T0 k� MC��G�&�1D"3Q	E1 4#Q ��O    ������HB�O�B�Ϻ	#�Io�Y|'�	���Em=����ǩ	/�3� T0 k� M_��c�&�1D"3Q	E1 4#Q ��O    ������PB�W�B�׺	'�Is�Y|'�	���Em?����ϩ	�3� T0 k� Mk��o�&�1D"3Q	E1 4#Q ��O    ������XB�_�E�ߺ	+�Is�Y|'�	���EmA����ө	�3� T0 k� -w��{�&�1D"3Q	E1 4#Q ��O    ������\B�g�E��	3�Is�Y|'�	|��EmD����۩	�3� T0 k� -�����&�1D"3Q	E1 4#Q ��O    ������dB�o�E��	7�Is�Y|'�	|��EmF�����	�3� T0 k� -�����&�1D"3Q	E1 4#Q  ��O    ������tB���E���?�Iw�Y|'�	|��E�K������#�3� T0 k� -�����&�1D"3Q	E1 4#Q# ��O    ������xB���E���C�Iw�Y|'�	|��E�M�������'�3� T0 k� ������&�1D"3Q	E1 4#Q$ ��O    ������B���E���K�Iw�Y|'�L��E�O������/�3� T0 k� ������&�1D"3Q	E1 4#Q% ��O    ������B͛�E���O�Iw�Y|'�L��E�R������3�3� T0 k� ������&�1D"3Q	E1 4#Q& ��O    ������ Bͣ�E�'��S�Iw�Y|'�L��E�T������7�3� T0 k� ������&�1D"3Q	E1 4#Q' ��O    ������ Bͫ�E�3��W�I{�Y|'�L��E�V������?�3� T0 k� ������&�1D"3Q	E1 4#Q( ��O    ������!Bͷ�E�;��_�I{�Y|'�L��E�Y����#��C�3� T0 k� ������&�1D"3Q	E1 4#Q) ��O    �������!BͿ�E�C��c�I{�Y|'�<��F[����+��K�3� T0 k� ����&�1D"3Q	E1 4#Q) ��O    �������!B�ǠE�O��g�I{�Y|'�<��F]����3�O�3� T0 k� .���&�1D"3Q	E1 4#Q* ��O    �������"B�ϠE�W��k�E�{�Y|'�<��F`����;�W�3� T0 k� .��#�&�1D"3Q	E1 4#Q+ ��O    �������#B�ߠE~k��w�E��Y|'�<��Fd����K�c�3� T0 k� .7��;�&�1D"3Q	E1 4#Q- ��O    �������#B��E~s��{�E��Y|'�<��Ff����S�g�3� T0 k� .C��G�&�1D"3Q	E1 4#Q. ��O    �������$B��E~{���E���Y|'�<��Fi����[�o�3� T0 k� �S��W�&�1D"3Q	E1 4#Q. ��O    �������$B���E~�����E���Y|'�<��Fk����c�s�3� T0 k� �_��c�&�1D"3Q	E1 4#Q/ ��O    �������%B��E~�����E���Y|+�<��Fm����k�{�3� T0 k� �k��o�&�1D"3Q	E1 4#Q0 ��O    �������%B��E~���� E���Y|+�<��Fp����s��3� T0 k� �t �x &�1D"3Q	E1 4#Q0 ��O    �������%B��E~��͐E���Y|+�,��Fr���{���3� T0 k� ����&�1D"3Q	E1 4#Q1 ��O    �������&B��E~��͔E���Y|+�,��Ft��߃���3� T0 k� ����&�1D"3Q	E1 4#Q2 ��O    ������&B�#�E~��͘B���Y|+�,��E�w��ߋ���3� T0 k� ����&�1D"3Q	E1 4#Q2 ��O    ������&B�+�E~��͜B���Y|+�,��E�y��ߓ���3� T0 k� ����&�1D"3Q	E1 4#Q3 ��    ������'B�7�E~��͜B���Y|+�,��E�{��ߛ���3� T0 k� .���&�1D"3Q	E1 4#Q3 ��    ������((B�G�En��ͤB���Y|+�,�E���߫���3� T0 k� .�	��	&�1D"3Q	E1 4#Q4 ��    ����� 0(B�O�En��ͨE���Y|+�,�E� ����߳����3� T0 k� .�
��
&�1D"3Q	E1 4#Q5 ��    ���   8(B�W�En��ͨ	E���Y|/�,�E�$����������3� T0 k� .���&�1D"3Q	E1 4#Q5 ��    ���  @)B�_�En��ͬ
E���Y|/�,�E�(�����é���3� T0 k� ����&�1D"3Q	E1 4#Q6 ��    ���  H)B�g�En��ͰE���Y|/�,�E�(�����˩���3� T0 k� � �&�1D"3Q	E1 4#Q6 ��    ���  P)B�s�En��ͰE���Y|/��
E�,����ө���3� T0 k� ��&�1D"3Q	E1 4#Q6 ��    ���  X*B�{�E���ݴE���Y|/��E�0����۩���3� T0 k� �� &�1D"3Q	E1 4#Q7 ��    ���  \*B���E���ݴDܻ�Y|/��E�4~��������3� T0 k� �(�,&�1D"3Q	E1 4#Q7 ��    ���  d*B���E���ݴDܿ�Y|/��E�8~����� ��3� T0 k� �4�8&�1D"3Q	E1 4#Q7 ��    ���  l+B���E��ݸD���Y|/��E�<}����� ��3� T0 k� �@�D&�1D"3Q	E1 4#Q7 ��    ���  t+B���E��ݸD���Y|/��E�@|������ ��3� T0 k� /P�T&�1D"3Q	E1 4#Q8 ��    ���   |+B���E��ݸD���Y|/��E�H|������ ��3� T0 k� /\�`&�1D"3Q	E1 4#Q8 ��    ��� # �,B���E���E���Y|/��E�L{����� �3� T0 k� /h�l&�1D"3Q	E1 4#Q8 ��    ��� & �,B���E���E���Y|/��B�Pz�˿�� �3� T0 k� /t�x&�1D"3Q	E1 4#Q8 ��    ��� ) �,B���E�#��E���Y|/��B�Ty�Ͼ�� �3� T0 k� /���&�1D"3Q	E1 4#Q8 ��    ��� , �-B�ǢE�'��E���Y|/��B�Xx�Ӿ�� �3� T0 k� ����&�1D"3Q	E1 4#Q8 ��    ��� 0 �-B�ϢE�+��E���Y|/���B�`w�ӽ�'� �3� T0 k� ����&�1D"3Q	E1 4#Q8 ��    ��� 3 �-B�ףF3��E���Y|/���B�dv�׽�/��#�3� T0 k� ����&�1D"3Q	E1 4#Q8 ��    ��� 6 �-B�ߣF7��E|��Y|, �� B�hv�ۼ�7��+�3� T0 k� �� �� &�1D"3Q	E1 4#Q8 ��    ��� 9 �.B��F;��E|��Y|, ��!B�pu�߼�?��3�3� T0 k� ��"��"&�1D"3Q	E1 4#Q8 ��    ��� < �.B��FC��E|��Y|, ��"B�ts���G��7�3� T0 k� ��#��#&�1D"3Q	E1 4#Q8 ��    ��� @ �.B���FG��E|��Y|, ��#B�xr���O��?�3� T0 k� ��$��$&�1D"3Q	E1 4#Q8 ��    ��� C �/B��FO��E}�Y|, ��$B��q���W��G�3� T0 k� /�&��&&�1D"3Q	E1 4#Q8 ��    ��� F �/B��FS��I��Y|, ��%B��p���_��O�3� T0 k� /�'��'&�1D"3Q	E1 4#Q8 ��    ��� I �/B��F[�� I��Y|, ��&B��o���g��S�3� T0 k�   (�(&�1D"3Q	E1 4#Q8 ��    ��� L �/B��F_��!I��Y|, ��'C�n����o��[�3� T0 k�  *�*&�1D"3Q	E1 4#Q8 ��    ��� P �0B�'�D�g��"I��Y|, ��(C�m����w��c�3� T0 k�  +� +&�1D"3Q	E1 4#Q8 ��    ��� S �0B�/�D�k��#I��Y|, ��)C�k������k�3� T0 k� �(,�,,&�1D"3Q	E1 4#Q6 ��    ��� V �0B�7�D�s��$I��Y|, ��*C�j������s�3� T0 k� �4-�8-&�1D"3Q	E1 4#Q6 ��    ��� Y �0B�?�D�w�m�%I��Y|, ��+C�i�� ���w�3� T0 k� �@/�D/&�1D"3Q	E1 4#Q6 ��    ��� \ �1B�G�D��m�&I��Y|, ��+C�h�� ����3� T0 k� �P0�T0&�1D"3Q	E1 4#Q5 ��    ��� ` �1B�O�D߀m�'I�#�Y|, ��,C�f�� �����3�T0 k� �\1�`1&�1D"3Q	E1 4#Q5 ��    ��� c �1B�W�D߈m�(I�#�Y|, ��,C�e�� �����3�T0 k� �h3�l3&�1D"3Q	E1 4#Q5 ��    ��� f �1B�c�Dߌm�)I�'�Y|, ��-E�c�� �����3�T0 k� �t4�x4&�1D"3Q	E1 4#Q4 ��    ��� i  1B�k�Dߔ}�*I�'�Y|, � -E�b�'� �����3�T0 k�  �5��5&�1D"3Q	E1 4#Q4 ��    ��� l 2B�s�Dߘ	}�,I�+�Y|, �.E�a�+� �����3�T0 k�  �7��7&�1D"3Q	E1 4#Q3 ��    �   p 2B�{�F�}�-I�+�Y|, �.E�`�3� ï���3�T0 k�  �8��8&�1D"3Q	E1 4#Q3 ��    �  s 2B߃�F�}�.I�/�Y|, �.E�^�7� ˰���3�T0 k�  �9��9&�1D"3Q	E1 4#Q3 ��    �  v 2Bߋ�F�}�/I�/�Y|, �.E�]�?� Ӱ���3�T0 k�  �;��;&�1D"3Q	E1 4#Q2 ��    �  y 3Bߓ�F�}�1I�/�Y|, �/E�\�G� ۱@��3�T0 k� ��<��<&�1D"3Q	E1 4#Q1 ��    �  } 3Bߟ�F�}�2I�3�Y|, �$/E�[�K��@��3�T0 k� ��=��=&�1D"3Q	E1 4#Q1 ��    �  �  3Bߧ�F���3I�3�Y|, �(/E Y�S��@��3�T0 k� ��?��?&�1D"3Q	E1 4#Q0 ��    �  � $3B߯�F���5I�3�Y|, �0/EX�[��@��3�T0 k� ��@��@&�1D"3Q	E1 4#Q0 ��    �  � ,3B߷�F���6I�3�Y|, �4/B�W�_���@��3�T0 k� ��A��A&�1D"3Q	E1 4#Q/ ��    �  � 03B߿�F���8I�3�Y|, �</B�V�g�� ���3�T0 k� �B�B&�1D"3Q	E1 4#Q. ��    � 	 � 44B�ǤE����9I�3�Y|, �D/B� U�o�� ���3�T0 k� �D�D&�1D"3Q	E1 4#Q. ��    � 
 � 84B�ϤE����;I�3�Y|, �H/B�(T�w�� ���3�T0 k� !E� E&�1D"3Q	E1 4#Q- ��    �  � <4B�ۤE����<I�3�Y|, �P.B�0S��� ���3�T0 k� !(F�,F&�1D"3Q	E1 4#Q, ��    �  � @4B��E��!��>A�3�Y|, �X.B�8Q���� ���3�T0 k� !4H�8H&�1D"3Q	E1 4#Q+ ��    �  � D4B��E��#��?A�3�Y|, �\.B�@P���'� ���3�T0 k� !DI�HI&�1D"3Q	E1 4#Q* ��    �  � H5B��B��$��AA�3�Y|, �d.B�HO���/� ��3�T0 k� !PJ�TJ&�1D"3Q	E1 4#Q* ��    �  � H5B���B� &��BA�3�Y|, �l-B�PN���!3� ��3�T0 k� �\L�`L&�1D"3Q	E1 4#Q) ��    �  � L5B��B�(�DA�3�Y|, �p-B�XM���!;� ��3�T0 k� �hM�lM&�1D"3Q	E1 4#Q( ��    �  � P5B��B�)�EA�3�Y|, �x,B�dL���!C� ��3�T0 k� �tN�xN&�1D"3Q	E1 4#Q' ��    �  � T5E��B�+�GA�3�Y|, ��,B�lK���!K� ��3�T0 k� ��P��P&�1D"3Q	E1 4#Q& ��    �  � X5E��B�-�HA�3�Y|, ��+B�tJ���!S� ��3�T0 k� ��Q��Q&�1D"3Q	E1 4#Q% ��    �  � \6E�'�B�$.�JA�3�Y|, ��+B�|J���![� �'�3�T0 k� ��R��R&�1D"3Q	E1 4#Q$ ��    �  � `6E�/�B�,0�KBM3�Y|, ��*B��I�Ǳ!_� �+�3�T0 k� ��T��T&�1D"3Q	E1 4#Q# ��    �  � d6E�7�B�41|LBM3�Y|, ��*B��Hϱ!g� �/��T0 k� !�U��U&�1D"3Q	E1 4#Q" ��    �  � d6E�?�B�<3xNBM3�Y|, ��)B��Gױ!o� �3��T0 k� !�V��V&�1D"3Q	E1 4#Q! �� 	   �  � h6E�K�B�D4tOBM3�Y|, ��(B��F߲!w� �;��T0 k� !�W��W&�1D"3Q	E1 4#Q  �� 	   �  � l6E�S�B�L6tPBM3�Y|, ��(B��E�!� �?��	T0 k� !�Y��Y&�1D"3Q	E1 4#Q �� 	   �  � p6E�[�B�T7pRBM3�Y|, ��'B��D��� �C��	T0 k� !�Z��Z&�1D"3Q	E1 4#Q �� 	   �  � t7E�c�B�\8lSBM3�Y|, ��'B��C���� �G��
T0 k� ��[��[&�1D"3Q	E1 4#Q �� 	   �  � t7B�k�B�d:dTBM3�Y|, ��&B��C���� �K��
T0 k� �]�]&�1D"3Q	E1 4#Q �� 	   �  � x7B�s�B�l;-`UBM3�Y|, ��&B��B��� �S��
T0 k� �^�^&�1D"3Q	E1 4#Q � 	   �  � |7B�{�B�t<-\W@3�Y|, ��%@�A��� �W��T0 k� �_� _&�1D"3Q	E1 4#Q � 	   �  � �7B���B�|>-XX@3�Y|, ��%@�@� a�� �[��T0 k� �(a�,a&�1D"3Q	E1 4#Q �� 	   �  � �7B���B��?-XY@3�Y|, ��$@�?#� a�� �_��T0 k� �4b�8b&�1D"3Q	E1 4#Q �� 	   �  � �7E��B��@-TZ@7�Y|,  �$@�?+� a�� �c��T0 k� �Dc�Hc&�1D"3Q	E1 4#Q �� 	   �  � �8E��B��BP[@7�Y|,  �#@�> 3� a�� �g��T0 k� "Pe�Te&�1D"3Q	E1 4#Q �� 	   �  � �8E��B��CL\B�7�Y|,  #@�= 7� a�� �k��T0 k� "\f�`f&�1D"3Q	E1 4#Q ��	   �  � �8E��B��DL]B�;�Y|,  "@ < ?� a�� �o��T0 k� "hg�lg&�1D"3Q	E1 4#Q �� 	   �  � �8E��B��EH^B�;�Y|,  "@< G� a�� �s��T0 k� "th�xh&�1D"3Q	E1 4#Q �� 	   �  � �8E��B��FH_B�;�Y|,  !@; O� a�� �w��T0 k� "�j��j&�1D"3Q	E1 4#Q �� 	   �  � �8EˠB��H�D`B�?�Y|,   !@: W� a�� �{��T0 k� ��k��k&�1D"3Q	E1 4#Q �� 	   �  � �8EӠB��I�DaB�?�Y|,  ( @ : _� a�� ���T0 k� ��l��l&�1D"3Q	E1 4#Q
 �� 	   �  � �8E�۟B��J�DbB�C�Y|,  0 @(9 c� a�� ����T0 k� ��n��n&�1D"3Q	E1 4#Q	 �� 	   �  � �9E��B��K�DcB�G�Y|,  8@,8 k� a�� ����T0 k� ��o��o&�1D"3Q	E1 4#Q �� 	   �  � �9E��B��L�@dB�G�Y|,  <@48 s� a�� ����T0 k� ��p��p&�1D"3Q	E1 4#Q �� 	   �  � �9E��B��M�@eB�K�Y|,  D@<7 w� a�� ����T0 k� ��r��r&�1D"3Q	E1 4#Q ��    �  � �9E���B��N�@fB�O�Y|,  L@D6 � a�� ����T0 k� ��s��s&�1D"3Q	E1 4#Q ��    �  � �9E��B��O�@gB�S�Y|,  P@H6 �� b� ����T0 k� "�t��t&�1D"3Q	E1 4#Q ��    �  � �9E��B�P�@hB�W�Y|,  X@P5 �� b� ����T0 k� "�v��v&�1D"3Q	E1 4#Q  ,�    �  � �9E��B�Q�@iB�[�Y|,  \@T4 �� b� ����T0 k� #w�w&�1D"3Q	E1 4#Q  ��    �  � �9E��B�R�@jB�_�Y|,  d@\4 �� b� ����T0 k� #x�x&�1D"3Q	E1 4#Q ��    �  � �9D�'�B� S�DkB�c�Y|,  h@d3 �� b� ����T0 k� #z� z&�1D"3Q	E1 4#Q ��    �  � �:D�/�B�(T�DlB�g�Y|,  p@h3 �� b� ����T0 k� �({�,{&�1D"3Q	E1 4#Q ��    �  � �:D�;�B�0U�DlB�k�Y|,  t@p2 �� b#� ����T0 k� �4|�8|&�1D"3Q	E1 4#Q ��    �  � �:D�C�B�<V�HmB�o�Y|,  |@t2 �� b'� ����T0 k� �D}�H}&�1D"3Q	E1 4#Q ��    �  � �:D�K�B�DW�HnB�s�Y|,  �@|1 �� b+� ����T0 k� �P�T&�1D"3Q	E1 4#Q ��    �  � �:D�S�B�LX�HoB�w�Y|,  �@�1 �� b/� ����T0 k� �\��`�&�1D"3Q	E1 4#Q ��    �  � �:D�[�B�TY�LpB��Y|,  �@�0 �� b7� ����T0 k� �h��l�&�1D"3Q	E1 4#Q ��    �  � �:D�c�B�`Z�LpB̓�Y|,  �@�/ Ǹ b;� ����T0 k� �t��x�&�1D"3Q	E1 4#Q *�    �  � �:D�k�B�hZ�PqB͇�Y|,  �@�/ ˹ b?� ����T0 k� �����&�1D"3Q	E1 4#Q ��    �  � �:D�s�B�p[�TrB͏�Y|,  �@�/ Ϲ bC� ����T0 k� �����&�1D"3Q	E1 4#Q ��    �  � �:D��B�x\�TsB͓�Y|,  �@�/ ׹ bG� ����T0 k� �����&�1D"3Q	E1 4#Q ��    �  � �;Dч�B��]�XsB͛�Y|,  �@�. ۹ bK� ����T0 k� �����&�1D"3Q	E1 4#Q ��    �  � �;DᏣB��^�\tB͟�a�,  �@�. ߹ bO� ���"c�T0 k� �����&�1D"3Q	E1 4#Q ��    �  � �;DᗣB��^�`uBͧ�a�,  �@�- � bS� ���"c�T0 k� ���ā&�1D"3Q	E1 4#Q ��    �  � �;D៤B��_�`vBͫ�a�,  �@�- � bW� ���"c�T0 k� �̀�Ѐ&�1D"3Q	E1 4#Q ��    �  � �;D᧤B��`�dvBݳ�a�,  �@�- � b[� ���"c�T0 k� �؀�܀&�1D"3Q	E1 4#Q ��    �  � �;DᯥB��a�hwBݷ�a�,  �@�, � b_� ���"c�T0 k� ����&�1D"3Q	E1 4#Q ��    �  � �;E���B��b�lxBݿ�a�,  �@�, �� bc� ���"c�T0 k� ����&�1D"3Q	E1 4#Q ��    �  � �;E���B��b�lxB���a�,  �@�+ �� bg� ���"c�T0 k� ��~� ~&�1D"3Q	E1 4#Q ��    �  � �;E�ǦB��c�pyB���a�,  �@�+ � bk� ���"c�T0 k� �|�|&�1D"3Q	E1 4#Q  ��   �  � �<E�ϧB��d�tyB���a�,  �@�* � bo� ���"c�T0 k� �{�{&�1D"3Q	E1 4#Q  ,�    �  � �<E�ۧB��d�tzB���a�,  �@�* � bs� ���"c�T0 k� �z� z&�1D"3Q	E1 4#Q  ��    �  � �<E��B��e�x{B���a�,  �@�) � bw� ���"c�T0 k� �$x�(x&�1D"3Q	E1 4#Q  ��    �  � �<E��B��f�|{B���Y|,  �@�) � b{� ����T0 k� �0w�4w&�1D"3Q	E1 4#Q  ��    �  � �<E��B��f�||B���Y|,  �@�) � b� ����T0 k� �8u�<u&�1D"3Q	E1 4#Q  ��    �  � �<Eq��B�g��}B���Y|,  �@�( � b�� ����T0 k� �@s�Ds&�1D"3Q	E1 4#Q  ��    �  � �<Er�B�h��}B��Y|,  �@�( � b�� ����T0 k� �Hq�Lq&�1D"3Q	E1 4#Q  ��    �  � �<Er�B�h��~B��Y|,  �@�' #� b�� ����T0 k� �Po�To&�1D"3Q	E1 4#Q  ��    �  � �<Er�E� i��~B��Y|,  �@�' '� b�� ����T0 k� �Xn�\n&�1D"3Q	E1 4#Q  ��    �  ���<Er�E�(j��B��Y|,  �@�' +� b�� ����T0 k� �\l�`l&�1D"3Q	E1 4#Q  ��    �  ���<D��E�4j��B��Y|,  �@�& /� b�� ����T0 k� �dj�hj&�1D"3Q	E1 4#Q  ��    �  ���=D�'�E�<k���B�'�Y|,  �@�& 3� b�� ����T0 k� �hh�lh&�1D"3Q	E1 4#Q  ��    �  ���=D�/�E�Hk���B�/�Y|,   @�& 7� b�� ����T0 k� �pf�tf&�1D"3Q	E1 4#Q  ��    �  ���=D�7�E�Pl��B�7�Y|,  @�% ;� b�� ����T0 k� �td�xd&�1D"3Q	E1 4#Q  ��    �  ���=D�?�E�Xm��B�?�a�,  @�% ?� b�� ���"C�T0 k� �xb�|b&�1D"3Q	E1 4#Q  ��    �  ���=D�C�E�dm��B�G�a�,  @�% ?� b�� ���"C�T0 k� �|`��`&�1D"3Q	E1 4#Q  ��    �  ���=D�K�E�ln��B�O�a�,  @�$ C� b�� ���"C�T0 k� ��^��^&�1D"3Q	E1 4#Q  ��    �  ���=D�S�E�tn��~B�W�a�,  @ $ G� b�� ���"C�T0 k� ��\��\&�1D"3Q	E1 4#Q  ��   �  ���=D�W�E��o��~B�_�a�,  @$ K� b�� ���"C�T0 k� ��Z��Z&�1D"3Q	E1 4#Q  ��    �  ���=D�_�E��o��~B�g�a�,  @# O� b�� ���"C�T0 k� ��X��X&�1D"3Q	E1 4#Q  ��    �  ���=D�c�E��p��~B�o�a�,  @# S� b�� ��"C�T0 k� ��V��V&�1D"3Q	E1 4#Q  ��    �  ���=D�k�E��p��}B�w�a�,  @# S� b�� ��"C�T0 k� ��T��T&�1D"3Q	E1 4#Q  ��    �  ���=D�s�E��p��}B��a�,   @" W� b�� ��"C�T0 k� ��R��R&�1D"3Q	E1 4#Q  ��    �  ���>D�w�E��p��}B���a�,  $@" [� b�� ��"C�T0 k� ��P��P&�1D"3Q	E1 4#Q  ��    �  ���>D��E��q��}B���a�,  (@" _� b�� ��"C�T0 k� ��N��N&�1D"3Q	E1 4#Q  ��    �  ���>D���E��q��}B���Y|,  ,@! _� b�� ���T0 k� ��L��L&�1D"3Q	E1 4#Q  ��    �  ���>D���E��q��|B���Y|,  ,@! c� b�� ���T0 k� ��J��J&�1D"3Q	E1 4#Q  ��    �  ���>D���E��q��|B���Y|,  0@ ! g� b�� ���T0 k� ��H��H&�1D"3Q	E1 4#Q  ��    �  ���>D���E��q��|B���Y|,  4@ ! k� b�� ���T0 k� ��F��F&�1D"3Q	E1 4#Q  ��    �  ���>D���E��q��|Bη�Y|,  4@$  k� b�� ���T0 k� ��D��D&�1D"3Q	E1 4#Q  ��    �  ���>D���E��q��|Bο�Y|,  8@(  o� b�� ���T0 k� ��B��B&�1D"3Q	E1 4#Q  ��    �  �� >D���E��q��{B���Y|,  <@(  s� b�� ���T0 k� ��@��@&�1D"3Q	E1 4#Q  ��    �  �� >D���E�q��{B���Y|,  <@,  s� b�� ���T0 k� ��>��>&�1D"3Q	E1 4#Q  ��    �  �� >D���E�p��{B���Y|,  @@0 w� b�� ���T0 k� ��<��<&�1D"3Q	E1 4#Q  ��    �  �� >D���E�p��{K���Y|,  D@0 {� b�� ���T0 k� ��;��;&�1D"3Q	E1 4#Q  ��    �  ��>D���E� p��{K���Y|,  D@4 {� b�� ���T0 k� ��9��9&�1D"3Q	E1 4#Q  ��    �  ��>D���E�(o��zK���Y|,  H@8 � b�� ���T0 k� ��7��7&�1D"3Q	E1 4#Q  ��    �  ��?D���E�0o��zK���Y|,  L@8 �� b�� ���T0 k� ��5��5&�1D"3Q	E1 4#Q  ��    �  ��?D���E�<n��zK���Y|,  L@< �� b�� ���T0 k� ��3��3&�1D"3Q	E1 4#Q  ��    �  ��?D���E�Dm��zK���Y|,  P@< �� b�� ���T0 k� ��2��2&�1D"3Q	E1 4#Q  ��    �  ��?D���E�Lm��zK��Y|,  P@@ �� b�� ���T0 k� ��0��0&�1D"3Q	E1 4#Q  ��    �  ��?D���E�Tl��zK��Y|,  T@@ �� b�� �#��T0 k� ��.��.&�1D"3Q	E1 4#Q  ��    �  ��?D���E�\k��yK��Y|,  X@D �� b�� �#��T0 k� ��,��,&�1D"3Q	E1 4#Q  ��    �  ��?D���E�`k��yK��Y|,  X@H �� b�� �#��T0 k� ��*��*&�1D"3Q	E1 4#Q  ��    �  ��?D���E�hj��yK��Y|,  \@H �� b�� �'��T0 k� ��)��)&�1D"3Q	E1 4#Q  ��    �  ��?D���E�pi��yK�#�Y|,  \@L �� b�� �'��T0 k� ��'��'&�1D"3Q	E1 4#Q  ��    �  ��?D���E�th��yK�+�Y|,  `@L �� b�� �'��T0 k� ��%��%&�1D"3Q	E1 4#Q  ��    �  ��?D���E�|g��yK�/�Y|,  `@P �� b�� �'��T0 k� ��#��#&�1D"3Q	E1 4#Q  ��    �  ��?D���EÄf��yK�7�Y|,  d@P �� b�� �+��T0 k� ��"��"&�1D"3Q	E1 4#Q  ��    �  ��?D���EÈe��xK�;�Y|,  d@T �� b�� �+��T0 k� �� �� &�1D"3Q	E1 4#Q  ��    �  ��?D���EÌd��xK�C�Y|,  h@T �� b�� �+��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��?D���EÔc��xK�G�Y|,  h@X �� b�� �/��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��?D���EØb��xK�K�Y|,  l@X �� b�� �/��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��?D���EÜa��xK�S�Y|,  l@\ �� b�� �/��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��?D���EӠ`��xK�W�Y|,  p@\ �� b�� �/��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@D���EӤ_��xK�[�Y|,  p@` �� b�� �3��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@D���EӨ^��xK�_�Y|,  t@` �� b�� �3��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@D��EӬ]��wK�g�Y|,  t@` �� c� �3��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@D��EӰ\��wK�k�Y|,  x@d �� c� �3��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@D��L�[��wK�o�Y|,  x@d �� c� �7��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@D��L�Z��wK�s�Y|,  x@h �� c  �7��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@D��L�Y��wK�s�Y|,  x@h �� c �7��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@D��L�Y��wK�w�Y|,  x@l �� c �7��T0 k� ��	��	&�1D"3Q	E1 4#Q  ��    �  ��@MS�L�X��wK�{�Y|,  |@l �� c �7��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@MS�L�W��wK��Y|,  |@l �� c �;��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@MS�L�V��vK���Y|,  �@p �� c �;��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@MS�L�U��vK���Y|,  �@p �� c �;��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@MS�L�T��vK���Y|,  �@p �� c �;��T0 k� ����&�1D"3Q	E1 4#Q  ��    �  ��@MS�L�S��vK���Y|,  �@t �� c	 �?��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��@MS#�L#�S� vK���Y|,  �@t �� c
 �?��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  � @MS'�L#�R�vK���Y|,  �@x �� c �?��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  � @MS'�L#�Q�vK���Y|,  �@x �� c �?��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  �  @MS+�L#�P�vK���Y|,  �@x �� c �?��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  �  @Mc+�L#�O�vK���Y|,  �@| �� c �C��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  �  @Mc/�L#�O�vK���Y|,  �@| �� c �C��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  �  @Mc/�L#�N�vK���Y|,  �@| �� c �C��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  �  @Mc3�L#�M� uK���Y|,  �@� �� c �C��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  �  @Mc4 L#�L�$uK���Y|,  �@� �� c �C��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  �  AMc4L#�L�(uK���Y|,  �@� �� c �G��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  � $AMc8L#�K�,uK���Y|,  �@� �� c  �G��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  � $AMc8L#�J�0uK���Y|,  �@� �� c  �G��T0 k� ������&�1D"3Q	E1 4#Q  ��    �  � $AMc<L$ J�4uK���Y|,  �@� �� c  �G�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  � $AMS<L$ I�8uK���Y|,  �@� �� c  �G�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  � $AMS@L$H�<uK���Y|,  �@� �� c$ �G�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  � $AMS@L$H�@uK���Y|,  �@� �� c$ �K�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  � $AMSDL$G�DuK���Y|,  �@� �� c$ �K�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��$AMSDL$F�HuK���Y|,  �@� �� c( �K�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��(AMSH	L$F�LuK���Y|,  �@� �� c( �K�� T0 k� ������&�1D"3Q	E1 4#Q  ��   �  ��(AMSH	L$E�PtK���Y|,  �@� �� c( �K�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��(AMSL
L$E�TtK���Y|,  �@� �� c( �K�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��(AMSLL$D�XtK���Y|,  �@� �� c, �K�� T0 k� ������&�1D"3Q	E1 4#Q  ��   �  ��(AD�PL$D�XtB���Y|,  �@� �� c, �O�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��(AD�PL$C�\tB���Y|,  �@� �� c, �O�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��(AD�PL$B�`tB���Y|,  �@� �� c, �O�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��(AD�TL$ B�dtB���Y|,  �@� �� c0 �O�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��(AD�TL$ A�htB���Y|,  �@� �� c0  �O�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��(AMSXL$$A�ltE���Y|,  �@� �� c0! �O�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��,AMSXL$$@�ltE���Y|,  �@� �� c0! �O�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  ��,AMS\L$(@�ptE���Y|,  �@� �� c4" �S�� T0 k� ������&�1D"3Q	E1 4#Q  ��    �  �                                                                                                                                                                            � � �  �  �  d A�  �K����   �      � \��%� ]�(p(o �  �� C`u   �       � ��     C_e �j      l           c  Z �           `�    ���   0
&


          |+  S S	     � ���     |�? �t    �^�k   	          Z �         �pb      ���  (
 
           i^�  S S	     �b     i2� �=`    ���             Z �         >�b     ��� 0	
           q��   + \	      fY     q�� 9�    �� �               Z �           ���    ���   H	$
          ��  � �
	   / _0=     �� ^�    !             6 Z �          �  &  ���  03 
            �0 ��	      C�3      �0�3           	                ����                 ���    P		 5              ��   T     W��O�     ����>�                            �          
@     ��@   (
	           ı  `       k 4S�     �� 4A�    W                     �          �      ��@   
	          ���  
     :    ��� +>       �                   ��           �@     ��@   8	 

          Hn�          � �Dn     H@M �Jh    ���              �         	 �      ��@   0
3
         ���        � �Y9    ��  �Pd     	 �                 � �         
       ��H   H


          #�� ��
     � ��     #�� ��     <                        ���l                ��@    		 5 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                         ����  ��        �     ��� o    �5��                    x                j  �   ��   �                         ��    ��        �      ��             "                                                �                           � �  _��� 4  � � ���   	 
              
    J�  ��D       �$ �e� �$ f� �D g  �d g  Є g@ Ф g` :� ``� ;D  a� ;� a� ;� b ���J ����X � AD �t� BD  u� B� v  � p�  p� � �t� � u� �d u� 
�< V� 
�| W  
�\ W  
�\ W� 
� W� 
�\ X  �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ���� ����� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��� �  ���4  ������  
�fD
��L���"����D"� �  " `   J jF��    "�j "���
��
���     �j��  
  �
� �  �  
� ��    ��     ��  �    C    ��     �       ����  ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �3&      ��&T ��        � �T ���        �        ��        �        ��        �    ��    ������'        ��                         T�) , 	 ��                                     �                 ����	            ������&��    � 2���2             18 Denis Savard e                                                                                   2  2     �C
2�BK/ �: K7 �B K8 �J K9 �2 K: �* K; �	c� �! 	c� �
J�OJ�_ J�G � J�P �K< �KL K4 � K= �c�$ �c�4 � c� �
c� � � c� � �	� � �	� � �� � �� �,"� �, "� �� � 
� � � *'{ � *'{ � *){ �"
� � #"L rD  " zz%*� � �&"�	 � '"� �(�	 �)
� �  "H r`  "J �S  "J �.-
� � � ."H rK  "J �^0") z^  "P �^  " zB3" zJ  "M �`  "S �G 6"M �_  "S � �8Bs ~ �9Bq � � :B� ~ � ;B� � v<Bo �.  "Q v  "C v �  *S                                                                                                                                                                                                                         x� P         �    @ 
        �     b P E e  ��         
            ������������������������������������� ���������	�
���������                                                                                          ��    �a�� ��������������������������������������������������������   �4, K   $@1�@A�A���j�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                2   ' '     �  ��J     \T                              ������������������������������������������������������                                                                                                                                           ����  ��                                             ������������������������� � ������������ ���������������  �� ������������� �������� ��������������� ��������������������������������������������������������������� ���������������� ����� ������������������������ ��  ������� �������                                   i    %    �� 
ĳJ      V�  	                           ������������������������������������������������������                                                                                                                                             ����  �  �                                           ��� ��� ��� �������������� �����������������  ������ �������� ��   ���������� ���������������������������  ��� ����� ���������  ������ �� ���� ������ � ��������� ����  ���  ����� ������������  ��� ��������������� �� �������                                                                                                                                                                                                                                                                   
                                                           �              


             �  }�         ���          N     6�                                                            ���^  6�      ,�����������������������������������������������������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � ��� �e�                                                                                                                                                                                                                                                                                      )n)n1n  
$              k      m                        l      m                                                                                                                                                                                                                                                                                                                                                                                                          > �  >�  J�  @�  -#�  EZm^  �N V����<����f���<��� �̎�o�̞������R�                 x � :�O        $   �   &  QW  �   �                    �                                                                                                                                                                                                                                                                                                                                        K K            -             !��                                                                                                                                                                                                                            Z   	�� �� Ѱ�      �� 4      ������������������������� � ������������ ���������������  �� ������������� �������� ��������������� ��������������������������������������������������������������� ���������������� ����� ������������������������ ��  ������� ���������� ��� ��� �������������� �����������������  ������ �������� ��   ���������� ���������������������������  ��� ����� ���������  ������ �� ���� ������ � ��������� ����  ���  ����� ������������  ��� ��������������� �� �������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     7   #   7   � ��                       4     �  ����������'      ��     T�      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ��    �� � �� �� �z � � �N ^$     �(        ��  �1   �    >�� ��  � ��   p �� �� �z   p���� �$ ^h  ��   p  � L��      +           �� �     ��   ��     �� A �� �� �z A ��  �� ��  O �� ��  �� ��  �� �� e� �� �� �z e� �$ �$ ^$         ��f&T  ��& T      �  ��   g���        f ^�         ��f       1      ��%����2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                                                  U  T   T   T     T UDUDDUDDDDDDDDDDDDDDDP   E�  DU� DDU�DDDUDDDDDDDDDDDD                UP  E�  E   E                                           ���U�UTD�DDDDDDTDD TDD   �   U_ DEU�DDDUDDDDD��DZT�DDDDDDDDDDDDTDDDDDDDDUTU�����DDDDDDDDDDDEDDDEDDDDTUTU�Ԫ���Z_   P   � �U�UTDUDDDDUTD�DT��D        U_��DEU_DDD_DDDPDDE�DDE  �DD DD DD �DD �UD  �U       DZTDEDDDDE�DDE�DDE�TDDT�DE�TE���DDTU�ZD���������DDTDD��ZT�T���ZTDDE��D��T�T��DUTTT��Z��TQTDDUTD�DDDTDDD�DDDDDDE�DD_TDE�DD_ DDP DDP DD_ DU_ U�  �                                       TE�DDD�UUU                    ���DDDUUUTD  D  D  D  D  U��D�TDDDDEUUDP  DP  DP  DP  UP  TDE�DDDPUUU_                                                    wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwtwwwCwwt1wwCwt1wC�t1��C1����������""""���������������!���""!����,���ww��7����������������wwwwwwwwwwwwwwwwwwww7wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwws��w1wt1�wC�t1��s��s��s������"$��Gw�!������������L���q��"r��������!�����!ww�r�w�ww!�wwrwwwwwwqwwwrwwww�7ww�ww�ww��7w��w���G��'!wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " ""  "!  " ! " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ ""   "! " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                            " ""   "" !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �              "   "   "�  �                        �   " ��.�  ��                   �                        ��"� �"� ����                  �  ".��".� ��                        ���          ���������������������  ��  ��  ��  �   �    �          �         �                                                                                              	�  �� �� ���ܙܽɪ�͚�����͙ͼ̨��̄DC"�D32�C33�333�33P330X̽ 
�� ˪  "   ""/"""�����vv ��p ��  ��  ̽  ˸  ɚ  ��  ؛  -�� .ܰ .��  �"  �   .   "�                   � �  ��            Z   Z   Z   Z  Z  �� �� �� "� "" "" ""/ ����   �   � .�". �" ����                    �� ��������p��r`     �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����         "� "     �  �   �   �         �     �                                                                                                                                                                                     	�  �� �� ���ܙܽɪ�͚�����͙ͼ̨��̄DC"�D32�C33�333�33P330X̽ 
�� ˪  "   ""/"""�����vv ��p ��  ��  ̽  ˸  ɚ  ��  ؛  -�� .ܰ .��  �"  �   .   "�                   � �  ��            Z   Z   Z   Z  Z  �� �� �� "� "" "" ""/ ����   �   � .�". �" ����                    �� ��������p��r`                �   ��  �ڛ�}ک�"   "   "  �� ��                   �".��".���                                ".  ".  ���   ��                                 � "�"  �    � � �                                                                                                                                                           ̙ �ɪ���˭�̻� �� �   ""  ""  .         �� ̻ �� ��w �rb �wg���z�����ٙ�����ˍ�ݙ8����DD��3D��33L�3� �3+ ��" �" ""  ".  �  �   �                        �T  �U  �D  +�� ��� 
�  �"" �"" ��"/��� ��� �  ��               �   �   �   �   �   �   �@      �    �  �   �""��""����         �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����            �   �   �   D   E�  U�  UO                         "  "  "      � "�"  �    � � �   �   "  "     "   "   �                                                                                                              �  �  �  �� ݚ� }�Ȫ��˙������˼� ��  ��  ��  ��  ��  I� H� �E X�T X�S T�D �[ ˻  ˸  ��  
� �,"��"" "  �" �  ""� �� ˻ �˻ ��ݪ��کɨ��ˀ�̽ ��� ��  ̽  ̻  ̻  ˉ  ��  �D  DC  C3  #;  ;�� �� ��  �� "�  "  �"/ / ����� ��  �      �   �          �  �  "     "  "  "   "�  �  �   �   
                            �          �   �          �                    �   �".� .�    ���.�                         �     �                                                                                                                                                                                          �  �  �  �  w  �  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �          �  .   �� ��     �  ��  �                         �� ��  �� �� ��� �           �   � �                   �         �  "� "  �  ��                                                                                                                                        �� ���
�������˽������̽�]��+I۲"T�""T32.T33>@4C CDT �E@ ��  ʐ  �       "   "�� � ��� �wp �&  �vz �w� �����˻���˰�̰� ��  ��  ��� � �+ �+ �  .   "�   �   �   �    � ��  �                     �  �˰ ���                 ".  ".  ���           U   U  U  U  	T  ,� ,� "  " "  ��  �            �"  �                        .   .   �                                           �    ���� �              .  ". ""  "    � ���                                                                                                                                                                                             �  ��� ��� }�� wݪ �� 	�� �� �ͼ ��� ��� ̘� �ͻ +���"�8"8  8� �� �U��EU��3 ̻�"̰""�" ��" �"                             �   ��� �˹��˚���ڍ�̽���ͽ��ͽ���ݼ��л�� ��D �UT EUT UU0 C3  2"  ""  -�  ��  ��  �   � ��"/ �" � ���    �        �   �   �"  "�  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                    ".  ".  ���                   ���                                      ���                          ����                  �   �� �       �  �  "�  "   "                                           �� �˨}��'ݪvw� w
�  
�  
�  �  �  "" �" " �  �                             ��        �   ��  ��� ��̰���˻�̻��̸̽��ۘ̚ɩ�D
��E˴EU�$PX"$ �"" �"" ɢ" 
��  �  "" """/����                             ��                                �                   �""��""�����    �  �  �           ���    �   �   E0  T4  S4@ 34@ CK� ��  ɫ  "̰�" �/ ���� ���                  �".��".  ���    �                    ".  ".  ���                   ���                                                                                                                                                                                                 	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                       ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �       �  �  �  �               ���                                                                                                                                                                                                           �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��r`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   �". ". ����                 �� �̽���ݪ۽w�}�&��vv���p��� ���  +"  "" ���������                   �                        ��"� �"� ����                            ".  ".  ���   ��                                 � "�"  �    � � �                            ����                  �   �� �       �  �  "�  "   "                                                             �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫒒 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          .� ".� "/� /�  �                         �   �                    �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                   2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD l � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=GwDGwqwDDwtwwww3333DDDD  � �!�aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( """"����������A��I��I X � �!�aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx""""�����A�DA�I��I� w � �!�aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""��������I���I���I���I��� � � �!�aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(MAMAMMMM�M�M����3333DDDD L  . M + , N    O P Q R S S S T S S S T S S 0 Z S ST S S ST S S SRQPO(( (N(,(+(M(.LD�����MD��M����3333DDDD  7  N 5 U V W X Y S S [ S S S _ S S S _ S S \ ] S S_ S S S_ S S S[ S SY(X(W(V(U(5(N((7���4���4���4���4���4���43334DDDD  `  V    a b c S S f g h i j i i i j i i ^ d i ij i i ij ihgf S Scb(a(((V((`""""wwwwqqqqwGwGGG 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
""""wwwwwwqqDAwG w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw������������������333DDD w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xwwM��M��D��M����������3333DDDD + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+DD��D�M��D����3333DDDD � W  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ������ ���((W(�""""������DH�H� � a � l � � � � � �������� � �� � � � � � ���	����� � � �� �������l(�(a(�""""�������H�H��D �  � y � � � � � � � � � � � � � � � �� ��������� � � � � � � � � ������y(�(�""""��������H��H��H��H� = l �  � � � � � � � � � � ��� � � � � �������� � � � ��� � � � ������((�l(=DD������L��DL����3333DDDD    �  � � � � � � � � � ������ � � � � � ���� � � � ������ � � �����((�(( L�A�AAD��DL�����3333DDDD x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���4���4���4L��4L��4���43334DDDD w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww""""���������M�MMM  � w w � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �����ww�(""""�������A��AA �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((���������������333DDD ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`I��I����������������3333DDDD M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M��A���I��I���I�����3333DDDD � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""������������������������ � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(�""""������D�D��� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5""""������������������������ x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�xwqwwqwwwwwqwwwDwwww3333DDDD w � � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxwwqqwwwDDwtGwwww3333DDDD � � � i i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+www4www4www4www4www4www43334DDDD W � � u u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(�""""wwwwwwqwwwqwqwq a � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�""""wwwwwwwDwGwA  � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(��A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDDC
2�BK/ �: K7 �B K8 �J K9 �2 K: �* K; �	c� �! 	c� �
J�OJ�_ J�G � J�P �K< �KL K4 � K= �c�$ �c�4 � c� �
c� � � c� � �	� � �	� � �� � �� �,"� �, "� �� � 
� � � *'{ � *'{ � *){ �"
� � #"L rD  " zz%*� � �&"�	 � '"� �(�	 �)
� �  "H r`  "J �S  "J �.-
� � � ."H rK  "J �^0") z^  "P �^  " zB3" zJ  "M �`  "S �G 6"M �_  "S � �8Bs ~ �9Bq � � :B� ~ � ;B� � v<Bo �.  "Q v  "C v �  *S3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ����>�L�L�T�\��=�L�S�H�U�U�L��������>��<���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���""""������A�D��I��""""�������D����� ��$��/�L�U�P�Z��=�H�]�H�Y�K���������>��<���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �8�>�7������A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �>��<��� ��""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II�""""������D""""������IADD���I""""��������D��""""�������I��I�I�I�""""�������A�D�II�I""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            